
module CONV_DW01_add_0 ( A, B, CI, SUM, CO );
  input [43:0] A;
  input [43:0] B;
  output [43:0] SUM;
  input CI;
  output CO;
  wire   \A[0] , n1, n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14,
         n15, n16, n17, n18, n19, n20, n21, n22, n23, n24, n25;
  wire   [43:1] carry;
  assign SUM[15] = A[15];
  assign SUM[14] = A[14];
  assign SUM[13] = A[13];
  assign SUM[12] = A[12];
  assign SUM[11] = A[11];
  assign SUM[10] = A[10];
  assign SUM[9] = A[9];
  assign SUM[8] = A[8];
  assign SUM[7] = A[7];
  assign SUM[6] = A[6];
  assign SUM[5] = A[5];
  assign SUM[4] = A[4];
  assign SUM[3] = A[3];
  assign SUM[2] = A[2];
  assign SUM[1] = A[1];
  assign \A[0]  = A[0];
  assign SUM[0] = \A[0] ;

  ADDFXL U1_23 ( .A(A[23]), .B(B[23]), .CI(n2), .CO(carry[24]), .S(SUM[23]) );
  ADDFXL U1_29 ( .A(A[29]), .B(B[29]), .CI(carry[29]), .CO(carry[30]), .S(
        SUM[29]) );
  ADDFXL U1_32 ( .A(A[32]), .B(B[32]), .CI(carry[32]), .CO(carry[33]), .S(
        SUM[32]) );
  ADDFXL U1_33 ( .A(A[33]), .B(B[33]), .CI(carry[33]), .CO(carry[34]), .S(
        SUM[33]) );
  ADDFXL U1_34 ( .A(A[34]), .B(B[34]), .CI(carry[34]), .CO(carry[35]), .S(
        SUM[34]) );
  ADDFXL U1_30 ( .A(A[30]), .B(B[30]), .CI(carry[30]), .CO(carry[31]), .S(
        SUM[30]) );
  ADDFXL U1_35 ( .A(A[35]), .B(B[35]), .CI(carry[35]), .CO(carry[36]), .S(
        SUM[35]) );
  ADDFHX2 U1_24 ( .A(A[24]), .B(B[24]), .CI(carry[24]), .CO(carry[25]), .S(
        SUM[24]) );
  CLKAND2X8 U1 ( .A(A[42]), .B(n23), .Y(n24) );
  NAND2X6 U2 ( .A(A[31]), .B(n4), .Y(n25) );
  BUFX8 U3 ( .A(carry[31]), .Y(n4) );
  NAND2X2 U4 ( .A(A[41]), .B(n10), .Y(n11) );
  INVX1 U5 ( .A(n22), .Y(n10) );
  CLKAND2X12 U6 ( .A(A[26]), .B(carry[26]), .Y(n17) );
  OR2X8 U7 ( .A(A[25]), .B(carry[25]), .Y(carry[26]) );
  BUFX4 U8 ( .A(carry[36]), .Y(n3) );
  NAND2X2 U9 ( .A(A[18]), .B(n1), .Y(n7) );
  CLKAND2X12 U10 ( .A(A[17]), .B(n14), .Y(n1) );
  XOR2X4 U11 ( .A(A[43]), .B(n24), .Y(SUM[43]) );
  CLKAND2X12 U12 ( .A(A[19]), .B(carry[19]), .Y(n15) );
  NAND3X4 U13 ( .A(n6), .B(n7), .C(n8), .Y(carry[19]) );
  CLKAND2X12 U14 ( .A(A[22]), .B(n13), .Y(n2) );
  NAND2X4 U15 ( .A(n11), .B(n12), .Y(SUM[41]) );
  AND2X2 U16 ( .A(A[37]), .B(n18), .Y(n19) );
  AND2X2 U17 ( .A(A[39]), .B(n20), .Y(n21) );
  AND2X2 U18 ( .A(A[21]), .B(carry[21]), .Y(n13) );
  OR2X2 U19 ( .A(A[20]), .B(n15), .Y(carry[21]) );
  AND2X2 U20 ( .A(A[36]), .B(n3), .Y(n18) );
  XOR2X1 U21 ( .A(A[42]), .B(n23), .Y(SUM[42]) );
  OR2X8 U22 ( .A(A[28]), .B(n16), .Y(carry[29]) );
  INVX4 U23 ( .A(n25), .Y(carry[32]) );
  XOR2X1 U24 ( .A(A[36]), .B(n3), .Y(SUM[36]) );
  CLKAND2X12 U25 ( .A(B[16]), .B(A[16]), .Y(n14) );
  XOR2XL U26 ( .A(B[18]), .B(A[18]), .Y(n5) );
  XOR2XL U27 ( .A(n1), .B(n5), .Y(SUM[18]) );
  NAND2X1 U28 ( .A(B[18]), .B(n1), .Y(n6) );
  NAND2XL U29 ( .A(A[18]), .B(B[18]), .Y(n8) );
  NAND2XL U30 ( .A(n9), .B(n22), .Y(n12) );
  CLKINVX1 U31 ( .A(A[41]), .Y(n9) );
  CLKAND2X12 U32 ( .A(A[40]), .B(n21), .Y(n22) );
  AND2X4 U33 ( .A(A[41]), .B(n22), .Y(n23) );
  XOR2XL U34 ( .A(A[40]), .B(n21), .Y(SUM[40]) );
  XOR2XL U35 ( .A(A[39]), .B(n20), .Y(SUM[39]) );
  XOR2XL U36 ( .A(A[38]), .B(n19), .Y(SUM[38]) );
  XOR2XL U37 ( .A(A[37]), .B(n18), .Y(SUM[37]) );
  XOR2XL U38 ( .A(A[31]), .B(n4), .Y(SUM[31]) );
  XOR2XL U39 ( .A(A[27]), .B(n17), .Y(SUM[27]) );
  XOR2XL U40 ( .A(A[26]), .B(carry[26]), .Y(SUM[26]) );
  XNOR2XL U41 ( .A(A[28]), .B(n16), .Y(SUM[28]) );
  XNOR2XL U42 ( .A(A[25]), .B(carry[25]), .Y(SUM[25]) );
  XOR2XL U43 ( .A(A[22]), .B(n13), .Y(SUM[22]) );
  XOR2XL U44 ( .A(A[19]), .B(carry[19]), .Y(SUM[19]) );
  XOR2XL U45 ( .A(A[21]), .B(carry[21]), .Y(SUM[21]) );
  XNOR2XL U46 ( .A(A[20]), .B(n15), .Y(SUM[20]) );
  XOR2XL U47 ( .A(A[17]), .B(n14), .Y(SUM[17]) );
  XOR2XL U48 ( .A(B[16]), .B(A[16]), .Y(SUM[16]) );
  AND2X2 U49 ( .A(A[27]), .B(n17), .Y(n16) );
  AND2X2 U50 ( .A(A[38]), .B(n19), .Y(n20) );
endmodule


module CONV_DW_cmp_0 ( A, B, TC, GE_LT, GE_GT_EQ, GE_LT_GT_LE, EQ_NE );
  input [19:0] A;
  input [19:0] B;
  input TC, GE_LT, GE_GT_EQ;
  output GE_LT_GT_LE, EQ_NE;
  wire   n119, n120, n121, n122, n123, n124, n125, n126, n127, n128, n129,
         n130, n131, n132, n133, n134, n135, n136, n137, n138, n139, n140,
         n141, n142, n143, n144, n145, n146, n147, n148, n149, n150, n151,
         n152, n153, n154, n155, n156, n157, n158, n159, n160, n161, n162,
         n163, n164, n165, n166, n167, n168, n169, n170, n171, n172, n173,
         n174, n175, n176, n177, n178;

  NOR2BX1 U55 ( .AN(B[2]), .B(A[2]), .Y(n173) );
  OAI222X4 U56 ( .A0(B[12]), .A1(n122), .B0(B[12]), .B1(n150), .C0(n122), .C1(
        n150), .Y(n149) );
  OAI222X2 U57 ( .A0(A[13]), .A1(n153), .B0(n153), .B1(n131), .C0(A[13]), .C1(
        n131), .Y(n152) );
  OAI222X4 U58 ( .A0(B[12]), .A1(n122), .B0(B[12]), .B1(n154), .C0(n154), .C1(
        n122), .Y(n153) );
  OAI22X4 U59 ( .A0(B[10]), .A1(n123), .B0(B[10]), .B1(n158), .Y(n157) );
  INVX2 U60 ( .A(n158), .Y(n124) );
  OAI222X4 U61 ( .A0(A[9]), .A1(n175), .B0(n175), .B1(n133), .C0(A[9]), .C1(
        n133), .Y(n158) );
  OAI222XL U62 ( .A0(B[17]), .A1(n120), .B0(B[17]), .B1(n178), .C0(n178), .C1(
        n120), .Y(n177) );
  OAI222XL U63 ( .A0(B[5]), .A1(n126), .B0(B[5]), .B1(n166), .C0(n126), .C1(
        n166), .Y(n165) );
  OAI222X1 U64 ( .A0(B[8]), .A1(n125), .B0(B[8]), .B1(n176), .C0(n176), .C1(
        n125), .Y(n175) );
  OAI222X1 U65 ( .A0(A[13]), .A1(n149), .B0(n131), .B1(n149), .C0(A[13]), .C1(
        n131), .Y(n148) );
  AOI2BB2X2 U66 ( .B0(n139), .B1(n140), .A0N(n137), .A1N(n119), .Y(n138) );
  OAI222X1 U67 ( .A0(B[14]), .A1(n121), .B0(B[14]), .B1(n148), .C0(n121), .C1(
        n148), .Y(n147) );
  NAND2BXL U68 ( .AN(B[7]), .B(A[7]), .Y(n176) );
  NOR2BXL U69 ( .AN(B[7]), .B(A[7]), .Y(n161) );
  INVX1 U70 ( .A(B[13]), .Y(n131) );
  INVX1 U71 ( .A(B[18]), .Y(n129) );
  OAI221XL U72 ( .A0(B[19]), .A1(n137), .B0(B[19]), .B1(n119), .C0(n138), .Y(
        GE_LT_GT_LE) );
  INVX1 U73 ( .A(A[8]), .Y(n125) );
  NAND2BXL U74 ( .AN(B[16]), .B(A[16]), .Y(n178) );
  NOR2BXL U75 ( .AN(B[16]), .B(A[16]), .Y(n143) );
  NAND2BXL U76 ( .AN(B[2]), .B(A[2]), .Y(n172) );
  AOI2BB1XL U77 ( .A0N(n136), .A1N(A[1]), .B0(B[0]), .Y(n174) );
  CLKINVX1 U78 ( .A(A[12]), .Y(n122) );
  CLKINVX1 U79 ( .A(n172), .Y(n128) );
  INVXL U80 ( .A(B[1]), .Y(n136) );
  CLKINVX1 U81 ( .A(A[5]), .Y(n126) );
  CLKINVX1 U82 ( .A(A[14]), .Y(n121) );
  CLKINVX1 U83 ( .A(A[17]), .Y(n120) );
  CLKINVX1 U84 ( .A(A[3]), .Y(n127) );
  INVXL U85 ( .A(B[11]), .Y(n132) );
  CLKINVX1 U86 ( .A(A[19]), .Y(n119) );
  CLKINVX1 U87 ( .A(A[10]), .Y(n123) );
  INVXL U88 ( .A(B[9]), .Y(n133) );
  INVXL U89 ( .A(B[4]), .Y(n135) );
  INVXL U90 ( .A(B[15]), .Y(n130) );
  INVXL U91 ( .A(B[6]), .Y(n134) );
  OAI21X1 U92 ( .A0(n144), .A1(n145), .B0(n146), .Y(n139) );
  AOI221X1 U93 ( .A0(A[10]), .A1(n124), .B0(n155), .B1(n156), .C0(n157), .Y(
        n144) );
  OAI222X1 U94 ( .A0(A[15]), .A1(n147), .B0(n130), .B1(n147), .C0(A[15]), .C1(
        n130), .Y(n146) );
  NAND2XL U95 ( .A(A[11]), .B(n132), .Y(n150) );
  OAI22XL U96 ( .A0(n119), .A1(n141), .B0(B[19]), .B1(n141), .Y(n140) );
  OAI21XL U97 ( .A0(A[18]), .A1(n129), .B0(n142), .Y(n141) );
  OAI22XL U98 ( .A0(n143), .A1(n120), .B0(B[17]), .B1(n143), .Y(n142) );
  OAI21XL U99 ( .A0(A[15]), .A1(n130), .B0(n151), .Y(n145) );
  OAI22XL U100 ( .A0(n152), .A1(n121), .B0(B[14]), .B1(n152), .Y(n151) );
  NOR2X1 U101 ( .A(n132), .B(A[11]), .Y(n154) );
  OAI22XL U102 ( .A0(n123), .A1(n159), .B0(B[10]), .B1(n159), .Y(n156) );
  OAI21XL U103 ( .A0(A[9]), .A1(n133), .B0(n160), .Y(n159) );
  OAI22XL U104 ( .A0(n161), .A1(n125), .B0(B[8]), .B1(n161), .Y(n160) );
  OAI21XL U105 ( .A0(n162), .A1(n163), .B0(n164), .Y(n155) );
  OAI222XL U106 ( .A0(A[6]), .A1(n165), .B0(n134), .B1(n165), .C0(A[6]), .C1(
        n134), .Y(n164) );
  NAND2X1 U107 ( .A(A[4]), .B(n135), .Y(n166) );
  OAI21XL U108 ( .A0(A[6]), .A1(n134), .B0(n167), .Y(n163) );
  OAI22XL U109 ( .A0(n168), .A1(n126), .B0(B[5]), .B1(n168), .Y(n167) );
  NOR2X1 U110 ( .A(n135), .B(A[4]), .Y(n168) );
  AOI221XL U111 ( .A0(A[3]), .A1(n128), .B0(n169), .B1(n170), .C0(n171), .Y(
        n162) );
  OAI22XL U112 ( .A0(B[3]), .A1(n127), .B0(B[3]), .B1(n172), .Y(n171) );
  OAI22XL U113 ( .A0(n173), .A1(n127), .B0(B[3]), .B1(n173), .Y(n170) );
  AO22X1 U114 ( .A0(n174), .A1(A[0]), .B0(A[1]), .B1(n136), .Y(n169) );
  OAI222XL U115 ( .A0(A[18]), .A1(n177), .B0(n177), .B1(n129), .C0(A[18]), 
        .C1(n129), .Y(n137) );
endmodule


module CONV_DW01_inc_1 ( A, SUM );
  input [20:0] A;
  output [20:0] SUM;

  wire   [20:2] carry;

  ADDHXL U1_1_19 ( .A(A[19]), .B(carry[19]), .CO(carry[20]), .S(SUM[19]) );
  ADDHXL U1_1_18 ( .A(A[18]), .B(carry[18]), .CO(carry[19]), .S(SUM[18]) );
  ADDHXL U1_1_17 ( .A(A[17]), .B(carry[17]), .CO(carry[18]), .S(SUM[17]) );
  ADDHXL U1_1_15 ( .A(A[15]), .B(carry[15]), .CO(carry[16]), .S(SUM[15]) );
  ADDHXL U1_1_14 ( .A(A[14]), .B(carry[14]), .CO(carry[15]), .S(SUM[14]) );
  ADDHXL U1_1_9 ( .A(A[9]), .B(carry[9]), .CO(carry[10]), .S(SUM[9]) );
  ADDHXL U1_1_8 ( .A(A[8]), .B(carry[8]), .CO(carry[9]), .S(SUM[8]) );
  ADDHXL U1_1_3 ( .A(A[3]), .B(carry[3]), .CO(carry[4]), .S(SUM[3]) );
  ADDHXL U1_1_16 ( .A(A[16]), .B(carry[16]), .CO(carry[17]), .S(SUM[16]) );
  ADDHXL U1_1_12 ( .A(A[12]), .B(carry[12]), .CO(carry[13]), .S(SUM[12]) );
  ADDHXL U1_1_11 ( .A(A[11]), .B(carry[11]), .CO(carry[12]), .S(SUM[11]) );
  ADDHXL U1_1_7 ( .A(A[7]), .B(carry[7]), .CO(carry[8]), .S(SUM[7]) );
  ADDHXL U1_1_6 ( .A(A[6]), .B(carry[6]), .CO(carry[7]), .S(SUM[6]) );
  ADDHXL U1_1_4 ( .A(A[4]), .B(carry[4]), .CO(carry[5]), .S(SUM[4]) );
  ADDHXL U1_1_2 ( .A(A[2]), .B(carry[2]), .CO(carry[3]), .S(SUM[2]) );
  ADDHXL U1_1_13 ( .A(A[13]), .B(carry[13]), .CO(carry[14]), .S(SUM[13]) );
  ADDHXL U1_1_10 ( .A(A[10]), .B(carry[10]), .CO(carry[11]), .S(SUM[10]) );
  ADDHXL U1_1_5 ( .A(A[5]), .B(carry[5]), .CO(carry[6]), .S(SUM[5]) );
  ADDHXL U1_1_1 ( .A(A[1]), .B(A[0]), .CO(carry[2]), .S(SUM[1]) );
  XOR2X1 U1 ( .A(carry[20]), .B(A[20]), .Y(SUM[20]) );
endmodule


module CONV_DW_mult_tc_2 ( a, b, product );
  input [19:0] a;
  input [19:0] b;
  output [39:0] product;
  wire   n1, n4, n5, n7, n9, n11, n12, n13, n15, n18, n19, n22, n23, n24, n25,
         n28, n29, n31, n34, n36, n37, n40, n41, n43, n46, n47, n48, n49, n51,
         n53, n55, n57, n58, n59, n61, n63, n64, n65, n67, n68, n69, n70, n71,
         n72, n73, n74, n75, n76, n77, n78, n79, n80, n81, n82, n83, n84, n85,
         n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96, n97, n98, n102,
         n103, n105, n107, n108, n109, n110, n111, n112, n113, n114, n115,
         n116, n117, n119, n121, n123, n124, n125, n126, n128, n130, n131,
         n132, n133, n134, n135, n136, n137, n138, n139, n140, n141, n142,
         n143, n144, n145, n146, n147, n150, n152, n153, n154, n155, n157,
         n159, n160, n162, n164, n165, n166, n167, n168, n169, n170, n171,
         n172, n173, n174, n176, n178, n180, n181, n182, n183, n184, n185,
         n188, n189, n190, n191, n193, n194, n195, n196, n197, n200, n201,
         n202, n203, n204, n205, n208, n209, n210, n211, n212, n213, n214,
         n215, n216, n217, n218, n219, n220, n222, n224, n225, n226, n227,
         n228, n229, n230, n231, n232, n233, n234, n235, n236, n237, n238,
         n239, n240, n241, n246, n247, n248, n249, n251, n252, n253, n254,
         n257, n258, n259, n260, n261, n262, n263, n264, n265, n266, n267,
         n268, n270, n271, n272, n273, n274, n275, n276, n277, n279, n280,
         n281, n282, n283, n286, n287, n289, n290, n291, n292, n293, n294,
         n296, n298, n299, n300, n301, n302, n303, n304, n305, n306, n307,
         n308, n309, n310, n311, n312, n313, n314, n315, n316, n318, n320,
         n321, n323, n325, n326, n327, n329, n331, n332, n333, n334, n335,
         n337, n338, n339, n341, n342, n343, n344, n345, n347, n349, n350,
         n351, n352, n353, n354, n356, n359, n364, n365, n366, n368, n370,
         n372, n374, n376, n377, n380, n381, n386, n388, n390, n391, n392,
         n393, n394, n395, n396, n397, n398, n399, n400, n401, n402, n403,
         n404, n405, n406, n407, n408, n409, n410, n411, n412, n413, n414,
         n415, n416, n417, n418, n419, n420, n421, n422, n423, n424, n425,
         n426, n427, n428, n429, n430, n431, n432, n433, n434, n435, n436,
         n437, n438, n439, n440, n441, n442, n443, n444, n445, n446, n447,
         n448, n449, n450, n451, n452, n453, n454, n455, n456, n457, n458,
         n459, n460, n461, n462, n463, n464, n465, n466, n467, n468, n469,
         n470, n471, n472, n473, n474, n475, n476, n477, n478, n479, n480,
         n481, n482, n483, n484, n485, n486, n487, n488, n489, n490, n491,
         n492, n493, n494, n495, n496, n497, n498, n499, n500, n501, n502,
         n503, n504, n505, n506, n507, n508, n509, n510, n511, n512, n513,
         n514, n515, n516, n517, n518, n519, n520, n521, n522, n523, n524,
         n525, n526, n527, n528, n529, n530, n531, n532, n533, n534, n535,
         n536, n537, n538, n539, n540, n541, n542, n543, n544, n545, n546,
         n547, n548, n549, n550, n551, n552, n553, n554, n555, n556, n557,
         n558, n559, n560, n561, n562, n563, n564, n565, n566, n567, n568,
         n569, n570, n571, n572, n573, n574, n575, n576, n577, n578, n579,
         n580, n581, n582, n583, n584, n585, n586, n587, n588, n589, n590,
         n591, n592, n593, n594, n595, n596, n597, n598, n599, n600, n601,
         n602, n603, n604, n605, n606, n607, n608, n609, n610, n611, n612,
         n613, n614, n615, n616, n617, n618, n619, n620, n621, n622, n623,
         n624, n625, n626, n627, n628, n629, n630, n631, n632, n633, n634,
         n635, n636, n637, n638, n639, n640, n641, n642, n643, n644, n645,
         n646, n647, n648, n649, n650, n651, n652, n653, n654, n655, n656,
         n657, n658, n659, n660, n661, n662, n663, n664, n665, n666, n667,
         n668, n669, n670, n671, n672, n673, n674, n675, n676, n677, n678,
         n679, n680, n681, n682, n683, n684, n685, n686, n687, n688, n689,
         n690, n691, n692, n693, n694, n695, n696, n697, n698, n699, n700,
         n701, n702, n703, n704, n705, n706, n707, n708, n709, n710, n711,
         n712, n713, n714, n715, n716, n717, n718, n719, n720, n721, n722,
         n723, n724, n725, n726, n727, n728, n729, n730, n731, n732, n733,
         n734, n735, n736, n737, n738, n739, n740, n741, n742, n743, n744,
         n745, n746, n747, n748, n749, n750, n751, n752, n753, n754, n755,
         n756, n757, n758, n759, n760, n761, n762, n763, n764, n765, n766,
         n767, n768, n769, n770, n771, n772, n773, n774, n775, n776, n777,
         n778, n779, n780, n781, n782, n783, n784, n785, n786, n787, n788,
         n789, n790, n791, n792, n793, n794, n795, n796, n797, n798, n799,
         n800, n801, n802, n803, n804, n805, n806, n807, n808, n809, n810,
         n811, n812, n813, n814, n815, n816, n817, n818, n819, n820, n821,
         n822, n823, n824, n825, n826, n827, n828, n829, n830, n831, n832,
         n833, n834, n835, n836, n837, n838, n839, n840, n841, n842, n843,
         n844, n845, n846, n847, n848, n849, n850, n851, n852, n853, n854,
         n855, n856, n857, n858, n859, n860, n861, n862, n863, n864, n865,
         n866, n867, n868, n869, n870, n871, n872, n873, n874, n875, n876,
         n877, n878, n879, n880, n881, n882, n883, n884, n885, n886, n887,
         n888, n889, n890, n891, n892, n893, n894, n895, n896, n897, n898,
         n899, n900, n901, n902, n903, n904, n905, n906, n907, n908, n909,
         n910, n911, n912, n913, n914, n915, n916, n917, n918, n919, n920,
         n921, n922, n923, n924, n925, n926, n927, n928, n929, n930, n931,
         n932, n933, n934, n935, n936, n937, n938, n939, n940, n941, n942,
         n943, n944, n945, n946, n947, n948, n949, n950, n951, n952, n953,
         n954, n955, n956, n957, n958, n959, n960, n961, n962, n963, n964,
         n965, n966, n967, n968, n969, n970, n971, n972, n973, n974, n975,
         n976, n977, n978, n979, n980, n981, n982, n983, n984, n985, n986,
         n987, n988, n989, n990, n991, n992, n993, n994, n995, n996, n997,
         n998, n999, n1001, n1002, n1003, n1004, n1005, n1006, n1007, n1008,
         n1009, n1010, n1011, n1012, n1013, n1014, n1015, n1016, n1017, n1018,
         n1019, n1020, n1021, n1022, n1023, n1024, n1025, n1026, n1027, n1028,
         n1029, n1030, n1032, n1033, n1034, n1036, \product[39] ,
         \product[38] , n1121, n1122, n1123, n1124, n1125, n1126, n1127, n1128,
         n1129, n1130, n1131, n1132, n1133, n1134, n1135, n1136, n1137, n1138,
         n1139, n1140, n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148,
         n1149, n1150, n1151, n1152, n1153, n1154, n1155, n1156, n1157, n1158,
         n1159, n1160, n1161, n1162, n1163, n1164, n1165, n1166, n1167, n1168,
         n1169, n1170, n1171, n1172, n1173, n1174, n1175, n1176, n1177, n1178,
         n1179, n1180, n1181, n1182, n1183, n1184, n1185, n1186, n1187, n1188,
         n1189, n1190, n1191, n1192, n1193, n1194, n1195, n1196, n1197, n1198,
         n1199, n1200, n1201, n1202, n1203, n1204, n1205, n1206, n1207, n1208,
         n1209, n1210, n1211, n1212, n1213, n1214, n1215, n1216, n1217, n1218,
         n1219, n1220, n1221, n1222, n1223, n1224, n1225, n1226, n1227, n1228,
         n1229, n1230, n1231, n1232, n1233, n1234, n1235, n1236, n1237, n1238,
         n1239, n1240, n1241, n1242, n1243, n1244, n1245, n1246, n1247;
  assign product[36] = \product[39] ;
  assign product[39] = \product[39] ;
  assign product[37] = \product[38] ;
  assign product[38] = \product[38] ;

  OAI21X4 U71 ( .A0(n166), .A1(n102), .B0(n103), .Y(n63) );
  XOR2X2 U948 ( .A(n131), .B(n67), .Y(product[32]) );
  INVX1 U949 ( .A(n314), .Y(n313) );
  XNOR2X2 U950 ( .A(n344), .B(n95), .Y(product[4]) );
  XOR2X4 U951 ( .A(n1222), .B(n1138), .Y(product[33]) );
  NAND2X2 U952 ( .A(n521), .B(n533), .Y(n267) );
  NOR2X2 U953 ( .A(n565), .B(n574), .Y(n289) );
  CMPR42X2 U954 ( .A(n791), .B(n759), .C(n577), .D(n568), .ICI(n573), .S(n565), 
        .ICO(n563), .CO(n564) );
  NOR2X4 U955 ( .A(n219), .B(n212), .Y(n210) );
  INVX1 U956 ( .A(n219), .Y(n217) );
  CLKBUFX6 U957 ( .A(n824), .Y(n1121) );
  NOR2X4 U958 ( .A(n208), .B(n184), .Y(n182) );
  CLKINVX3 U959 ( .A(n210), .Y(n208) );
  NAND2X2 U960 ( .A(n365), .B(n364), .Y(n184) );
  AOI21X2 U961 ( .A0(n1125), .A1(n262), .B0(n263), .Y(n261) );
  OAI21X1 U962 ( .A0(n272), .A1(n264), .B0(n267), .Y(n263) );
  OAI22X1 U963 ( .A0(n936), .A1(n18), .B0(n935), .B1(n15), .Y(n757) );
  OAI22XL U964 ( .A0(n935), .A1(n18), .B0(n934), .B1(n15), .Y(n756) );
  XNOR2X1 U965 ( .A(n989), .B(n13), .Y(n935) );
  XOR2X4 U966 ( .A(n299), .B(n87), .Y(product[12]) );
  BUFX8 U967 ( .A(n889), .Y(n1122) );
  XNOR2X1 U968 ( .A(n997), .B(n31), .Y(n889) );
  CMPR42X1 U969 ( .A(n638), .B(n410), .C(n414), .D(n652), .ICI(n411), .S(n408), 
        .ICO(n406), .CO(n407) );
  ADDFX2 U970 ( .A(n666), .B(n416), .CI(n681), .CO(n409), .S(n410) );
  NOR2X1 U971 ( .A(n803), .B(n632), .Y(n353) );
  NAND2X4 U972 ( .A(n803), .B(n632), .Y(n354) );
  OAI22X2 U973 ( .A0(n982), .A1(n5), .B0(n981), .B1(n4), .Y(n803) );
  NAND2XL U974 ( .A(n235), .B(n238), .Y(n78) );
  OAI21X1 U975 ( .A0(n230), .A1(n238), .B0(n231), .Y(n229) );
  NAND2X2 U976 ( .A(n472), .B(n482), .Y(n238) );
  XNOR2X1 U977 ( .A(n990), .B(n7), .Y(n954) );
  BUFX16 U978 ( .A(a[10]), .Y(n990) );
  XNOR2X4 U979 ( .A(n994), .B(n19), .Y(n922) );
  NAND2X1 U980 ( .A(n419), .B(n413), .Y(n164) );
  CMPR42X2 U981 ( .A(n667), .B(n639), .C(n415), .D(n422), .ICI(n418), .S(n413), 
        .ICO(n411), .CO(n412) );
  NOR2X2 U982 ( .A(n259), .B(n266), .Y(n257) );
  NOR2X2 U983 ( .A(n521), .B(n533), .Y(n266) );
  XNOR2X4 U984 ( .A(n239), .B(n78), .Y(product[21]) );
  OAI21X4 U985 ( .A0(n248), .A1(n252), .B0(n249), .Y(n247) );
  NAND2X2 U986 ( .A(n496), .B(n507), .Y(n252) );
  NAND2X6 U987 ( .A(n483), .B(n495), .Y(n249) );
  BUFX12 U988 ( .A(n932), .Y(n1205) );
  XNOR2X2 U989 ( .A(n986), .B(n13), .Y(n932) );
  NAND2X2 U990 ( .A(n442), .B(n451), .Y(n213) );
  ADDHX2 U991 ( .A(n801), .B(n631), .CO(n621), .S(n622) );
  OAI22X1 U992 ( .A0(n980), .A1(n5), .B0(n979), .B1(n4), .Y(n801) );
  NOR2BX1 U993 ( .AN(n61), .B(n9), .Y(n786) );
  CLKBUFX12 U994 ( .A(a[0]), .Y(n61) );
  XNOR2X4 U995 ( .A(n987), .B(n1), .Y(n969) );
  BUFX12 U996 ( .A(a[13]), .Y(n987) );
  OAI22X2 U997 ( .A0(n874), .A1(n41), .B0(n873), .B1(n40), .Y(n696) );
  OAI22X2 U998 ( .A0(n1126), .A1(n40), .B0(n873), .B1(n41), .Y(n695) );
  XNOR2X1 U999 ( .A(n999), .B(n37), .Y(n873) );
  CLKBUFX6 U1000 ( .A(n877), .Y(n1209) );
  BUFX8 U1001 ( .A(n907), .Y(n1206) );
  XNOR2X1 U1002 ( .A(n997), .B(n25), .Y(n907) );
  OAI22X1 U1003 ( .A0(n969), .A1(n5), .B0(n968), .B1(n4), .Y(n790) );
  OAI22X4 U1004 ( .A0(n967), .A1(n4), .B0(n968), .B1(n1020), .Y(n789) );
  NOR2X4 U1005 ( .A(n442), .B(n451), .Y(n212) );
  NAND2X4 U1006 ( .A(n188), .B(n1130), .Y(n173) );
  OR2X2 U1007 ( .A(n420), .B(n425), .Y(n1130) );
  CLKBUFX6 U1008 ( .A(n876), .Y(n1123) );
  NOR2X4 U1009 ( .A(n400), .B(n402), .Y(n138) );
  CMPR42X2 U1010 ( .A(n650), .B(n404), .C(n665), .D(n636), .ICI(n401), .S(n400), .ICO(n398), .CO(n399) );
  CMPR42X2 U1011 ( .A(n405), .B(n637), .C(n409), .D(n651), .ICI(n406), .S(n403), .ICO(n401), .CO(n402) );
  NOR2X2 U1012 ( .A(n403), .B(n407), .Y(n145) );
  OAI22X1 U1013 ( .A0(n965), .A1(n1029), .B0(n12), .B1(n1142), .Y(n631) );
  NAND2X4 U1014 ( .A(n246), .B(n228), .Y(n226) );
  AOI21X4 U1015 ( .A0(n247), .A1(n228), .B0(n229), .Y(n227) );
  NOR2X2 U1016 ( .A(n237), .B(n230), .Y(n228) );
  NAND2X2 U1017 ( .A(n217), .B(n220), .Y(n76) );
  OAI21X4 U1018 ( .A0(n212), .A1(n220), .B0(n213), .Y(n211) );
  NAND2X2 U1019 ( .A(n452), .B(n460), .Y(n220) );
  XNOR2X2 U1020 ( .A(n984), .B(n7), .Y(n948) );
  BUFX12 U1021 ( .A(a[16]), .Y(n984) );
  AO21X4 U1022 ( .A0(n257), .A1(n274), .B0(n258), .Y(n1243) );
  OAI21X1 U1023 ( .A0(n259), .A1(n267), .B0(n260), .Y(n258) );
  OAI22X1 U1024 ( .A0(n879), .A1(n36), .B0(n878), .B1(n34), .Y(n700) );
  XNOR2X2 U1025 ( .A(n986), .B(n31), .Y(n878) );
  NAND2X4 U1026 ( .A(n434), .B(n441), .Y(n202) );
  CMPR42X2 U1027 ( .A(n457), .B(n453), .C(n454), .D(n445), .ICI(n450), .S(n442), .ICO(n440), .CO(n441) );
  XNOR2X2 U1028 ( .A(n985), .B(n7), .Y(n949) );
  BUFX20 U1029 ( .A(a[15]), .Y(n985) );
  OAI22X2 U1030 ( .A0(n913), .A1(n22), .B0(n914), .B1(n24), .Y(n735) );
  XNOR2X2 U1031 ( .A(n986), .B(n19), .Y(n914) );
  OAI22X2 U1032 ( .A0(n983), .A1(n4), .B0(n5), .B1(n1173), .Y(n632) );
  NAND2BXL U1033 ( .AN(n61), .B(n1), .Y(n983) );
  XNOR2X2 U1034 ( .A(n986), .B(n1), .Y(n968) );
  OAI22X1 U1035 ( .A0(n980), .A1(n4), .B0(n981), .B1(n5), .Y(n802) );
  NAND2X4 U1036 ( .A(n1174), .B(n1175), .Y(n980) );
  BUFX8 U1037 ( .A(n842), .Y(n1124) );
  XNOR2X1 U1038 ( .A(n986), .B(n43), .Y(n842) );
  XOR2X4 U1039 ( .A(n1247), .B(n79), .Y(product[20]) );
  CLKINVX8 U1040 ( .A(n201), .Y(n365) );
  NOR2X6 U1041 ( .A(n173), .B(n201), .Y(n171) );
  NOR2X4 U1042 ( .A(n434), .B(n441), .Y(n201) );
  CMPR42X2 U1043 ( .A(n644), .B(n479), .C(n718), .D(n687), .ICI(n473), .S(n464), .ICO(n462), .CO(n463) );
  OAI22X1 U1044 ( .A0(n1203), .A1(n1016), .B0(n896), .B1(n28), .Y(n718) );
  NAND2X2 U1045 ( .A(n224), .B(n210), .Y(n204) );
  AOI21X2 U1046 ( .A0(n225), .A1(n210), .B0(n211), .Y(n205) );
  NAND2X4 U1047 ( .A(n210), .B(n171), .Y(n169) );
  NOR2X2 U1048 ( .A(n452), .B(n460), .Y(n219) );
  CMPR42X2 U1049 ( .A(n466), .B(n462), .C(n463), .D(n455), .ICI(n459), .S(n452), .ICO(n450), .CO(n451) );
  NOR2X6 U1050 ( .A(n433), .B(n426), .Y(n190) );
  CMPR42X2 U1051 ( .A(n684), .B(n443), .C(n437), .D(n444), .ICI(n440), .S(n434), .ICO(n432), .CO(n433) );
  NAND2X4 U1052 ( .A(n1214), .B(n1215), .Y(n896) );
  CLKAND2X3 U1053 ( .A(n257), .B(n273), .Y(n1242) );
  OAI22X2 U1054 ( .A0(n946), .A1(n1018), .B0(n945), .B1(n15), .Y(n767) );
  INVX12 U1055 ( .A(n63), .Y(\product[39] ) );
  OR2X2 U1056 ( .A(n885), .B(n1015), .Y(n1220) );
  INVX3 U1057 ( .A(n994), .Y(n1165) );
  NAND2X4 U1058 ( .A(n1147), .B(n1148), .Y(n814) );
  CLKBUFX3 U1059 ( .A(n1013), .Y(n47) );
  CLKBUFX4 U1060 ( .A(b[13]), .Y(n37) );
  CLKBUFX3 U1061 ( .A(n1014), .Y(n41) );
  BUFX2 U1062 ( .A(n1019), .Y(n12) );
  OAI22X1 U1063 ( .A0(n926), .A1(n23), .B0(n925), .B1(n1027), .Y(n747) );
  OAI22X1 U1064 ( .A0(n977), .A1(n5), .B0(n976), .B1(n4), .Y(n798) );
  OAI22X1 U1065 ( .A0(n978), .A1(n5), .B0(n977), .B1(n4), .Y(n799) );
  OAI22X2 U1066 ( .A0(n960), .A1(n11), .B0(n959), .B1(n9), .Y(n781) );
  OAI22X1 U1067 ( .A0(n975), .A1(n4), .B0(n976), .B1(n5), .Y(n797) );
  INVX1 U1068 ( .A(n320), .Y(n318) );
  NAND2X1 U1069 ( .A(n224), .B(n195), .Y(n193) );
  INVXL U1070 ( .A(n619), .Y(n1219) );
  INVX3 U1071 ( .A(n343), .Y(n341) );
  OR2X2 U1072 ( .A(n886), .B(n34), .Y(n1160) );
  OR2X1 U1073 ( .A(n885), .B(n34), .Y(n1216) );
  OR2X1 U1074 ( .A(n888), .B(n36), .Y(n1157) );
  BUFX8 U1075 ( .A(n940), .Y(n1207) );
  OAI22X1 U1076 ( .A0(n951), .A1(n12), .B0(n950), .B1(n1029), .Y(n772) );
  OAI22XL U1077 ( .A0(n836), .A1(n51), .B0(n837), .B1(n53), .Y(n662) );
  CMPR42X1 U1078 ( .A(n528), .B(n516), .C(n754), .D(n722), .ICI(n522), .S(n511), .ICO(n509), .CO(n510) );
  CMPR42X1 U1079 ( .A(n689), .B(n720), .C(n646), .D(n503), .ICI(n704), .S(n489), .ICO(n487), .CO(n488) );
  CMPR42X1 U1080 ( .A(n491), .B(n500), .C(n736), .D(n504), .ICI(n497), .S(n486), .ICO(n484), .CO(n485) );
  OAI22XL U1081 ( .A0(n846), .A1(n48), .B0(n845), .B1(n46), .Y(n670) );
  NAND2X1 U1082 ( .A(n1181), .B(n1182), .Y(n890) );
  CLKBUFX3 U1083 ( .A(n922), .Y(n1204) );
  CLKINVX1 U1084 ( .A(n190), .Y(n188) );
  CMPR42X1 U1085 ( .A(n539), .B(n527), .C(n536), .D(n524), .ICI(n532), .S(n521), .ICO(n519), .CO(n520) );
  CLKINVX1 U1086 ( .A(n416), .Y(n417) );
  CMPR42X1 U1087 ( .A(n658), .B(n686), .C(n701), .D(n672), .ICI(n458), .S(n455), .ICO(n453), .CO(n454) );
  OAI22XL U1088 ( .A0(n1208), .A1(n51), .B0(n832), .B1(n53), .Y(n658) );
  OAI22XL U1089 ( .A0(n849), .A1(n47), .B0(n848), .B1(n1023), .Y(n673) );
  OAI21X1 U1090 ( .A0(n275), .A1(n281), .B0(n276), .Y(n274) );
  NAND2X1 U1091 ( .A(n1168), .B(n1169), .Y(n1171) );
  CMPR42X1 U1092 ( .A(n680), .B(n695), .C(n790), .D(n569), .ICI(n758), .S(n559), .ICO(n557), .CO(n558) );
  CMPR42X1 U1093 ( .A(n726), .B(n710), .C(n742), .D(n774), .ICI(n571), .S(n562), .ICO(n560), .CO(n561) );
  CMPR42X1 U1094 ( .A(n729), .B(n627), .C(n588), .D(n592), .ICI(n777), .S(n586), .ICO(n584), .CO(n585) );
  OAI22XL U1095 ( .A0(n955), .A1(n1029), .B0(n956), .B1(n11), .Y(n777) );
  XOR2X1 U1096 ( .A(b[10]), .B(b[11]), .Y(n1005) );
  NAND2X1 U1097 ( .A(n1141), .B(n1142), .Y(n1144) );
  AOI21X1 U1098 ( .A0(n225), .A1(n195), .B0(n196), .Y(n194) );
  OR2X1 U1099 ( .A(n286), .B(n289), .Y(n1245) );
  OA21X2 U1100 ( .A0(n286), .A1(n290), .B0(n287), .Y(n1246) );
  OAI22XL U1101 ( .A0(n843), .A1(n46), .B0(n844), .B1(n48), .Y(n668) );
  CMPR42X1 U1102 ( .A(n467), .B(n477), .C(n474), .D(n464), .ICI(n470), .S(n461), .ICO(n459), .CO(n460) );
  NOR2X2 U1103 ( .A(n461), .B(n471), .Y(n230) );
  ADDFHX2 U1104 ( .A(n800), .B(n768), .CI(n784), .CO(n619), .S(n620) );
  OAI22XL U1105 ( .A0(n964), .A1(n11), .B0(n963), .B1(n9), .Y(n785) );
  NAND2X1 U1106 ( .A(n136), .B(n1131), .Y(n125) );
  NAND2X1 U1107 ( .A(n1129), .B(n1127), .Y(n154) );
  CLKINVX1 U1108 ( .A(n121), .Y(n119) );
  NAND2X1 U1109 ( .A(n123), .B(n1132), .Y(n116) );
  AOI21X2 U1110 ( .A0(n306), .A1(n314), .B0(n307), .Y(n305) );
  OAI22XL U1111 ( .A0(n973), .A1(n5), .B0(n972), .B1(n4), .Y(n794) );
  CLKINVX1 U1112 ( .A(n331), .Y(n329) );
  CMPR42X1 U1113 ( .A(n765), .B(n629), .C(n749), .D(n611), .ICI(n612), .S(n609), .ICO(n607), .CO(n608) );
  NAND2X1 U1114 ( .A(n1177), .B(n1178), .Y(n765) );
  CLKXOR2X2 U1115 ( .A(n277), .B(n83), .Y(product[16]) );
  XOR2X2 U1116 ( .A(n261), .B(n81), .Y(product[18]) );
  OR2X1 U1117 ( .A(n419), .B(n413), .Y(n1129) );
  OAI21XL U1118 ( .A0(n155), .A1(n134), .B0(n135), .Y(n133) );
  NOR2X1 U1119 ( .A(n597), .B(n603), .Y(n311) );
  NAND2X1 U1120 ( .A(n622), .B(n785), .Y(n349) );
  NAND2X1 U1121 ( .A(n1176), .B(n352), .Y(n350) );
  OR2X1 U1122 ( .A(n354), .B(n351), .Y(n1176) );
  NOR2X1 U1123 ( .A(n802), .B(n786), .Y(n351) );
  NOR2X1 U1124 ( .A(n392), .B(n391), .Y(n111) );
  NOR2X1 U1125 ( .A(n116), .B(n111), .Y(n109) );
  INVX1 U1126 ( .A(n303), .Y(n301) );
  CLKINVX1 U1127 ( .A(n305), .Y(n304) );
  NAND2X1 U1128 ( .A(n597), .B(n603), .Y(n312) );
  CLKXOR2X2 U1129 ( .A(n339), .B(n94), .Y(product[5]) );
  CLKINVX1 U1130 ( .A(n1218), .Y(n338) );
  NAND2XL U1131 ( .A(n365), .B(n202), .Y(n74) );
  INVX1 U1132 ( .A(n202), .Y(n200) );
  BUFX2 U1133 ( .A(n282), .Y(n1125) );
  INVX1 U1134 ( .A(n283), .Y(n282) );
  OA21X2 U1135 ( .A0(n253), .A1(n251), .B0(n252), .Y(n1247) );
  XNOR2X1 U1136 ( .A(n987), .B(n43), .Y(n843) );
  OAI22XL U1137 ( .A0(n843), .A1(n48), .B0(n1124), .B1(n46), .Y(n667) );
  OAI22X1 U1138 ( .A0(n841), .A1(n46), .B0(n1124), .B1(n48), .Y(n666) );
  OAI22XL U1139 ( .A0(n854), .A1(n1023), .B0(n855), .B1(n47), .Y(n678) );
  XNOR2X1 U1140 ( .A(n998), .B(n43), .Y(n854) );
  BUFX3 U1141 ( .A(n872), .Y(n1126) );
  OAI22X1 U1142 ( .A0(n858), .A1(n40), .B0(n859), .B1(n1014), .Y(n416) );
  BUFX20 U1143 ( .A(a[2]), .Y(n998) );
  INVX1 U1144 ( .A(n13), .Y(n1169) );
  OR2X2 U1145 ( .A(n412), .B(n408), .Y(n1127) );
  OR2X1 U1146 ( .A(n609), .B(n613), .Y(n1128) );
  CLKBUFX3 U1147 ( .A(b[5]), .Y(n13) );
  XNOR2X1 U1148 ( .A(n993), .B(n25), .Y(n903) );
  OAI22X1 U1149 ( .A0(n852), .A1(n47), .B0(n851), .B1(n1023), .Y(n675) );
  CLKBUFX3 U1150 ( .A(n1020), .Y(n5) );
  CLKBUFX3 U1151 ( .A(n1012), .Y(n53) );
  XNOR2X2 U1152 ( .A(b[6]), .B(b[5]), .Y(n1027) );
  NAND2X2 U1153 ( .A(n1008), .B(n1028), .Y(n1018) );
  NAND2X2 U1154 ( .A(n1005), .B(n1025), .Y(n1015) );
  OR2X1 U1155 ( .A(n399), .B(n395), .Y(n1131) );
  OR2X1 U1156 ( .A(n394), .B(n393), .Y(n1132) );
  OR2X1 U1157 ( .A(n622), .B(n785), .Y(n1133) );
  OR2X1 U1158 ( .A(n614), .B(n615), .Y(n1134) );
  INVXL U1159 ( .A(n155), .Y(n153) );
  INVX1 U1160 ( .A(n154), .Y(n152) );
  OR2X2 U1161 ( .A(n604), .B(n608), .Y(n1135) );
  OR2X2 U1162 ( .A(n575), .B(n582), .Y(n1136) );
  XNOR2X1 U1163 ( .A(n994), .B(n25), .Y(n904) );
  BUFX4 U1164 ( .A(b[9]), .Y(n25) );
  CLKBUFX4 U1165 ( .A(b[17]), .Y(n49) );
  CLKINVX1 U1166 ( .A(n7), .Y(n1142) );
  CLKBUFX3 U1167 ( .A(b[1]), .Y(n1) );
  BUFX4 U1168 ( .A(b[15]), .Y(n43) );
  CLKBUFX3 U1169 ( .A(b[11]), .Y(n31) );
  CLKBUFX3 U1170 ( .A(b[19]), .Y(n55) );
  OR2X1 U1171 ( .A(n633), .B(n390), .Y(n1137) );
  NAND2X2 U1172 ( .A(n1006), .B(n1026), .Y(n1016) );
  NAND2X1 U1173 ( .A(n1001), .B(n1021), .Y(n1011) );
  CLKBUFX3 U1174 ( .A(n1011), .Y(n59) );
  BUFX6 U1175 ( .A(a[12]), .Y(n988) );
  CLKINVX1 U1176 ( .A(n302), .Y(n300) );
  CLKINVX1 U1177 ( .A(n337), .Y(n335) );
  NOR2X1 U1178 ( .A(n275), .B(n280), .Y(n273) );
  NOR2X1 U1179 ( .A(n620), .B(n621), .Y(n342) );
  XNOR2X1 U1180 ( .A(n997), .B(n37), .Y(n871) );
  XNOR2X1 U1181 ( .A(n997), .B(n19), .Y(n925) );
  XNOR2X1 U1182 ( .A(n986), .B(n37), .Y(n860) );
  XNOR2X1 U1183 ( .A(n993), .B(n19), .Y(n921) );
  XNOR2X1 U1184 ( .A(n991), .B(n1), .Y(n973) );
  INVX3 U1185 ( .A(n227), .Y(n225) );
  XNOR2X1 U1186 ( .A(n995), .B(n55), .Y(n815) );
  OAI22X1 U1187 ( .A0(n893), .A1(n34), .B0(n36), .B1(n1180), .Y(n627) );
  NAND2X1 U1188 ( .A(n1143), .B(n1144), .Y(n961) );
  NOR2X2 U1189 ( .A(n472), .B(n482), .Y(n237) );
  XNOR2X2 U1190 ( .A(b[2]), .B(b[1]), .Y(n1029) );
  AND2X2 U1191 ( .A(n1132), .B(n121), .Y(n1138) );
  XNOR2X1 U1192 ( .A(n988), .B(n7), .Y(n952) );
  XNOR2X1 U1193 ( .A(n999), .B(n49), .Y(n837) );
  OAI22X1 U1194 ( .A0(n899), .A1(n1016), .B0(n898), .B1(n28), .Y(n720) );
  OAI22XL U1195 ( .A0(n918), .A1(n24), .B0(n917), .B1(n22), .Y(n739) );
  XNOR2X1 U1196 ( .A(n990), .B(n19), .Y(n918) );
  XNOR2X1 U1197 ( .A(n985), .B(n37), .Y(n859) );
  XNOR2X1 U1198 ( .A(n985), .B(n43), .Y(n841) );
  XNOR2X1 U1199 ( .A(n998), .B(n13), .Y(n944) );
  CMPR42X2 U1200 ( .A(n501), .B(n489), .C(n498), .D(n486), .ICI(n494), .S(n483), .ICO(n481), .CO(n482) );
  OR2X1 U1201 ( .A(n138), .B(n146), .Y(n1139) );
  NAND2X2 U1202 ( .A(n1139), .B(n139), .Y(n137) );
  AOI21X2 U1203 ( .A0(n137), .A1(n1131), .B0(n128), .Y(n126) );
  AND2X2 U1204 ( .A(n165), .B(n109), .Y(n1140) );
  NOR2X6 U1205 ( .A(n1140), .B(n110), .Y(n108) );
  OAI21X2 U1206 ( .A0(n117), .A1(n111), .B0(n112), .Y(n110) );
  NAND2X1 U1207 ( .A(n997), .B(n7), .Y(n1143) );
  INVX1 U1208 ( .A(n997), .Y(n1141) );
  NAND2X1 U1209 ( .A(n994), .B(n55), .Y(n1147) );
  NAND2X2 U1210 ( .A(n1145), .B(n1146), .Y(n1148) );
  INVX1 U1211 ( .A(n994), .Y(n1145) );
  CLKINVX1 U1212 ( .A(n55), .Y(n1146) );
  OR2X6 U1213 ( .A(n814), .B(n57), .Y(n1227) );
  NOR2X1 U1214 ( .A(n879), .B(n34), .Y(n1149) );
  NOR2X1 U1215 ( .A(n880), .B(n36), .Y(n1150) );
  OR2X1 U1216 ( .A(n1149), .B(n1150), .Y(n701) );
  NOR2X1 U1217 ( .A(n924), .B(n22), .Y(n1151) );
  NOR2X1 U1218 ( .A(n925), .B(n23), .Y(n1152) );
  OR2X4 U1219 ( .A(n1151), .B(n1152), .Y(n746) );
  OR2X1 U1220 ( .A(n921), .B(n23), .Y(n1153) );
  OR2X1 U1221 ( .A(n920), .B(n22), .Y(n1154) );
  NAND2X1 U1222 ( .A(n1153), .B(n1154), .Y(n742) );
  BUFX12 U1223 ( .A(a[5]), .Y(n995) );
  OR2X1 U1224 ( .A(n910), .B(n29), .Y(n1155) );
  OR2X1 U1225 ( .A(n909), .B(n28), .Y(n1156) );
  NAND2X2 U1226 ( .A(n1155), .B(n1156), .Y(n731) );
  OR2X4 U1227 ( .A(n887), .B(n34), .Y(n1158) );
  NAND2X2 U1228 ( .A(n1157), .B(n1158), .Y(n709) );
  OR2X2 U1229 ( .A(n887), .B(n1015), .Y(n1159) );
  NAND2X6 U1230 ( .A(n1159), .B(n1160), .Y(n708) );
  ADDFHX4 U1231 ( .A(n708), .B(n788), .CI(n693), .CO(n541), .S(n542) );
  OR2XL U1232 ( .A(n933), .B(n15), .Y(n1161) );
  OR2XL U1233 ( .A(n934), .B(n18), .Y(n1162) );
  NAND2X2 U1234 ( .A(n1161), .B(n1162), .Y(n755) );
  XNOR2X2 U1235 ( .A(n987), .B(n13), .Y(n933) );
  XNOR2X1 U1236 ( .A(n988), .B(n13), .Y(n934) );
  NOR2X1 U1237 ( .A(n957), .B(n11), .Y(n1163) );
  NOR2X1 U1238 ( .A(n956), .B(n9), .Y(n1164) );
  OR2X1 U1239 ( .A(n1163), .B(n1164), .Y(n778) );
  NAND2X2 U1240 ( .A(n994), .B(n13), .Y(n1166) );
  NAND2X6 U1241 ( .A(n1165), .B(n1169), .Y(n1167) );
  NAND2X6 U1242 ( .A(n1166), .B(n1167), .Y(n940) );
  NAND2XL U1243 ( .A(n61), .B(n13), .Y(n1170) );
  NAND2X2 U1244 ( .A(n1170), .B(n1171), .Y(n946) );
  INVXL U1245 ( .A(n61), .Y(n1168) );
  NAND2XL U1246 ( .A(n998), .B(n1), .Y(n1174) );
  NAND2X1 U1247 ( .A(n1172), .B(n1173), .Y(n1175) );
  INVXL U1248 ( .A(n998), .Y(n1172) );
  INVXL U1249 ( .A(n1), .Y(n1173) );
  OR2XL U1250 ( .A(n944), .B(n1018), .Y(n1177) );
  OR2X1 U1251 ( .A(n943), .B(n15), .Y(n1178) );
  NAND2XL U1252 ( .A(n998), .B(n31), .Y(n1181) );
  NAND2X1 U1253 ( .A(n1179), .B(n1180), .Y(n1182) );
  INVXL U1254 ( .A(n998), .Y(n1179) );
  INVXL U1255 ( .A(n31), .Y(n1180) );
  OAI22X1 U1256 ( .A0(n890), .A1(n34), .B0(n891), .B1(n1015), .Y(n712) );
  NOR2X1 U1257 ( .A(n864), .B(n41), .Y(n1183) );
  NOR2X1 U1258 ( .A(n863), .B(n40), .Y(n1184) );
  OR2X1 U1259 ( .A(n1183), .B(n1184), .Y(n686) );
  NOR2X1 U1260 ( .A(n906), .B(n29), .Y(n1185) );
  NOR2X1 U1261 ( .A(n905), .B(n28), .Y(n1186) );
  OR2X1 U1262 ( .A(n1185), .B(n1186), .Y(n727) );
  NAND2XL U1263 ( .A(n990), .B(n1), .Y(n1188) );
  NAND2X1 U1264 ( .A(n1187), .B(n1173), .Y(n1189) );
  NAND2X1 U1265 ( .A(n1188), .B(n1189), .Y(n972) );
  INVXL U1266 ( .A(n990), .Y(n1187) );
  OAI22XL U1267 ( .A0(n972), .A1(n5), .B0(n971), .B1(n4), .Y(n793) );
  OR2X1 U1268 ( .A(n313), .B(n311), .Y(n1190) );
  NAND2X2 U1269 ( .A(n1190), .B(n312), .Y(n310) );
  OR2X6 U1270 ( .A(n155), .B(n125), .Y(n1191) );
  NAND2X8 U1271 ( .A(n1191), .B(n126), .Y(n124) );
  NAND2XL U1272 ( .A(n988), .B(n43), .Y(n1193) );
  NAND2X1 U1273 ( .A(n1192), .B(n1033), .Y(n1194) );
  NAND2X1 U1274 ( .A(n1193), .B(n1194), .Y(n844) );
  INVXL U1275 ( .A(n988), .Y(n1192) );
  OAI22X1 U1276 ( .A0(n845), .A1(n48), .B0(n844), .B1(n46), .Y(n669) );
  NAND2XL U1277 ( .A(n998), .B(n19), .Y(n1197) );
  NAND2X1 U1278 ( .A(n1195), .B(n1196), .Y(n1198) );
  NAND2X2 U1279 ( .A(n1197), .B(n1198), .Y(n926) );
  INVXL U1280 ( .A(n998), .Y(n1195) );
  INVXL U1281 ( .A(n19), .Y(n1196) );
  CLKBUFX3 U1282 ( .A(b[7]), .Y(n19) );
  OAI22X1 U1283 ( .A0(n926), .A1(n1027), .B0(n927), .B1(n23), .Y(n748) );
  NAND2XL U1284 ( .A(n988), .B(n49), .Y(n1199) );
  NAND2X1 U1285 ( .A(n1192), .B(n1032), .Y(n1200) );
  NAND2X1 U1286 ( .A(n1199), .B(n1200), .Y(n826) );
  OAI22X1 U1287 ( .A0(n827), .A1(n53), .B0(n826), .B1(n51), .Y(n653) );
  OR2X4 U1288 ( .A(n941), .B(n1018), .Y(n1201) );
  OR2X1 U1289 ( .A(n1207), .B(n15), .Y(n1202) );
  NAND2X2 U1290 ( .A(n1201), .B(n1202), .Y(n762) );
  CMPR42X2 U1291 ( .A(n762), .B(n746), .C(n778), .D(n714), .ICI(n600), .S(n594), .ICO(n592), .CO(n593) );
  OA21X4 U1292 ( .A0(n253), .A1(n222), .B0(n227), .Y(n1228) );
  INVX6 U1293 ( .A(n254), .Y(n253) );
  NOR2X1 U1294 ( .A(n154), .B(n125), .Y(n123) );
  OA21X1 U1295 ( .A0(n253), .A1(n193), .B0(n194), .Y(n1237) );
  OAI22X2 U1296 ( .A0(n923), .A1(n23), .B0(n1204), .B1(n1027), .Y(n744) );
  OAI22X2 U1297 ( .A0(n924), .A1(n23), .B0(n923), .B1(n22), .Y(n745) );
  CMPR42X2 U1298 ( .A(n659), .B(n674), .C(n645), .D(n703), .ICI(n688), .S(n478), .ICO(n476), .CO(n477) );
  OAI22X1 U1299 ( .A0(n834), .A1(n53), .B0(n833), .B1(n51), .Y(n659) );
  OA21X4 U1300 ( .A0(n253), .A1(n180), .B0(n181), .Y(n1232) );
  NAND2XL U1301 ( .A(n224), .B(n182), .Y(n180) );
  ADDHX4 U1302 ( .A(n781), .B(n797), .CO(n610), .S(n611) );
  XNOR2X1 U1303 ( .A(n990), .B(n13), .Y(n936) );
  NOR2X2 U1304 ( .A(n248), .B(n251), .Y(n246) );
  NOR2X4 U1305 ( .A(n483), .B(n495), .Y(n248) );
  OAI22X1 U1306 ( .A0(n854), .A1(n47), .B0(n853), .B1(n46), .Y(n677) );
  XNOR2X1 U1307 ( .A(n993), .B(n55), .Y(n813) );
  OAI22X4 U1308 ( .A0(n869), .A1(n41), .B0(n868), .B1(n40), .Y(n691) );
  XNOR2X2 U1309 ( .A(n994), .B(n37), .Y(n868) );
  OAI22X1 U1310 ( .A0(n867), .A1(n41), .B0(n866), .B1(n1024), .Y(n689) );
  XNOR2X1 U1311 ( .A(n987), .B(n19), .Y(n915) );
  NOR2X6 U1312 ( .A(n950), .B(n12), .Y(n1231) );
  XNOR2X4 U1313 ( .A(n986), .B(n7), .Y(n950) );
  BUFX4 U1314 ( .A(n897), .Y(n1203) );
  OAI21X1 U1315 ( .A0(n253), .A1(n240), .B0(n241), .Y(n239) );
  CMPR42X2 U1316 ( .A(n717), .B(n468), .C(n733), .D(n643), .ICI(n465), .S(n458), .ICO(n456), .CO(n457) );
  OAI22X2 U1317 ( .A0(n833), .A1(n53), .B0(n832), .B1(n51), .Y(n468) );
  OAI22X1 U1318 ( .A0(n917), .A1(n24), .B0(n916), .B1(n22), .Y(n738) );
  OAI22X4 U1319 ( .A0(n870), .A1(n41), .B0(n869), .B1(n40), .Y(n692) );
  XNOR2X2 U1320 ( .A(n995), .B(n37), .Y(n869) );
  OAI22X1 U1321 ( .A0(n838), .A1(n53), .B0(n837), .B1(n51), .Y(n663) );
  XNOR2X1 U1322 ( .A(n995), .B(n31), .Y(n887) );
  OAI22X1 U1323 ( .A0(n1203), .A1(n28), .B0(n898), .B1(n1016), .Y(n719) );
  AOI21X1 U1324 ( .A0(n165), .A1(n132), .B0(n133), .Y(n131) );
  XNOR2X1 U1325 ( .A(n988), .B(n1), .Y(n970) );
  OAI21X1 U1326 ( .A0(n253), .A1(n204), .B0(n205), .Y(n203) );
  OA21X4 U1327 ( .A0(n291), .A1(n289), .B0(n290), .Y(n1240) );
  OAI22X1 U1328 ( .A0(n955), .A1(n12), .B0(n954), .B1(n9), .Y(n776) );
  XNOR2X1 U1329 ( .A(n991), .B(n7), .Y(n955) );
  OAI22X4 U1330 ( .A0(n931), .A1(n15), .B0(n1205), .B1(n18), .Y(n753) );
  OAI22X1 U1331 ( .A0(n933), .A1(n18), .B0(n1205), .B1(n15), .Y(n754) );
  XNOR2X1 U1332 ( .A(n995), .B(n13), .Y(n941) );
  AOI21X2 U1333 ( .A0(n211), .A1(n171), .B0(n172), .Y(n170) );
  NOR2X2 U1334 ( .A(n208), .B(n197), .Y(n195) );
  XNOR2X1 U1335 ( .A(n992), .B(n7), .Y(n956) );
  BUFX12 U1336 ( .A(a[8]), .Y(n992) );
  OAI21X1 U1337 ( .A0(n173), .A1(n202), .B0(n174), .Y(n172) );
  XNOR2X1 U1338 ( .A(n998), .B(n49), .Y(n836) );
  XNOR2X1 U1339 ( .A(n993), .B(n31), .Y(n885) );
  OAI22X1 U1340 ( .A0(n905), .A1(n29), .B0(n904), .B1(n28), .Y(n726) );
  OAI22X1 U1341 ( .A0(n859), .A1(n40), .B0(n860), .B1(n41), .Y(n682) );
  OAI22X1 U1342 ( .A0(n861), .A1(n41), .B0(n860), .B1(n40), .Y(n683) );
  XNOR2X4 U1343 ( .A(n310), .B(n89), .Y(product[10]) );
  AOI21X1 U1344 ( .A0(n200), .A1(n364), .B0(n189), .Y(n185) );
  BUFX12 U1345 ( .A(a[3]), .Y(n997) );
  OAI21X2 U1346 ( .A0(n227), .A1(n169), .B0(n170), .Y(n168) );
  XNOR2X1 U1347 ( .A(n994), .B(n49), .Y(n832) );
  XOR2X4 U1348 ( .A(n268), .B(n82), .Y(product[17]) );
  BUFX20 U1349 ( .A(a[7]), .Y(n993) );
  XNOR2X1 U1350 ( .A(n995), .B(n49), .Y(n833) );
  OAI22X1 U1351 ( .A0(n890), .A1(n1015), .B0(n1122), .B1(n34), .Y(n711) );
  OAI22X4 U1352 ( .A0(n1209), .A1(n34), .B0(n878), .B1(n36), .Y(n699) );
  XNOR2X1 U1353 ( .A(n165), .B(n71), .Y(product[28]) );
  ADDFHX4 U1354 ( .A(n752), .B(n493), .CI(n660), .CO(n490), .S(n491) );
  INVX3 U1355 ( .A(n492), .Y(n493) );
  AOI21X4 U1356 ( .A0(n1130), .A1(n189), .B0(n176), .Y(n174) );
  OAI21X1 U1357 ( .A0(n308), .A1(n312), .B0(n309), .Y(n307) );
  OAI22X1 U1358 ( .A0(n852), .A1(n46), .B0(n853), .B1(n47), .Y(n676) );
  ADDHX2 U1359 ( .A(n745), .B(n761), .CO(n587), .S(n588) );
  OAI21X1 U1360 ( .A0(n253), .A1(n233), .B0(n234), .Y(n232) );
  XNOR2X1 U1361 ( .A(n989), .B(n1), .Y(n971) );
  XNOR2X1 U1362 ( .A(n999), .B(n19), .Y(n927) );
  BUFX12 U1363 ( .A(a[1]), .Y(n999) );
  XNOR2X1 U1364 ( .A(n993), .B(n13), .Y(n939) );
  CMPR42X2 U1365 ( .A(n550), .B(n540), .C(n547), .D(n537), .ICI(n543), .S(n534), .ICO(n532), .CO(n533) );
  ADDFHX2 U1366 ( .A(n780), .B(n764), .CI(n796), .CO(n605), .S(n606) );
  OAI22X1 U1367 ( .A0(n959), .A1(n11), .B0(n958), .B1(n9), .Y(n780) );
  ADDFHX2 U1368 ( .A(n735), .B(n492), .CI(n751), .CO(n479), .S(n480) );
  BUFX3 U1369 ( .A(n831), .Y(n1208) );
  OAI22X1 U1370 ( .A0(n906), .A1(n28), .B0(n1206), .B1(n29), .Y(n728) );
  OAI22X1 U1371 ( .A0(n908), .A1(n29), .B0(n1206), .B1(n28), .Y(n729) );
  XOR2X4 U1372 ( .A(n140), .B(n68), .Y(product[31]) );
  OAI22X1 U1373 ( .A0(n978), .A1(n4), .B0(n979), .B1(n5), .Y(n800) );
  NOR2X4 U1374 ( .A(n508), .B(n520), .Y(n259) );
  XOR2X4 U1375 ( .A(n113), .B(n65), .Y(product[34]) );
  OAI22X1 U1376 ( .A0(n942), .A1(n15), .B0(n943), .B1(n1018), .Y(n764) );
  CMPR42X2 U1377 ( .A(n724), .B(n756), .C(n678), .D(n552), .ICI(n740), .S(n540), .ICO(n538), .CO(n539) );
  OAI22X1 U1378 ( .A0(n903), .A1(n29), .B0(n902), .B1(n28), .Y(n724) );
  OAI22X1 U1379 ( .A0(n975), .A1(n5), .B0(n974), .B1(n4), .Y(n796) );
  XNOR2X1 U1380 ( .A(n995), .B(n7), .Y(n959) );
  XOR2X4 U1381 ( .A(n160), .B(n70), .Y(product[29]) );
  OAI21X2 U1382 ( .A0(n253), .A1(n215), .B0(n216), .Y(n214) );
  OAI22X2 U1383 ( .A0(n951), .A1(n1029), .B0(n952), .B1(n12), .Y(n773) );
  XNOR2X1 U1384 ( .A(n987), .B(n7), .Y(n951) );
  OAI21X1 U1385 ( .A0(n209), .A1(n184), .B0(n185), .Y(n183) );
  CMPR42X2 U1386 ( .A(n624), .B(n541), .C(n531), .D(n538), .ICI(n535), .S(n527), .ICO(n525), .CO(n526) );
  OAI22X1 U1387 ( .A0(n839), .A1(n51), .B0(n53), .B1(n1032), .Y(n624) );
  XOR2X4 U1388 ( .A(n108), .B(n64), .Y(product[35]) );
  CMPR42X2 U1389 ( .A(n696), .B(n572), .C(n579), .D(n576), .ICI(n570), .S(n568), .ICO(n566), .CO(n567) );
  ADDHX1 U1390 ( .A(n727), .B(n743), .CO(n571), .S(n572) );
  CMPR42X2 U1391 ( .A(n725), .B(n694), .C(n553), .D(n679), .ICI(n741), .S(n551), .ICO(n549), .CO(n550) );
  OAI22X1 U1392 ( .A0(n903), .A1(n28), .B0(n904), .B1(n29), .Y(n725) );
  OAI22X1 U1393 ( .A0(n928), .A1(n23), .B0(n927), .B1(n1027), .Y(n749) );
  OAI21X1 U1394 ( .A0(n209), .A1(n197), .B0(n202), .Y(n196) );
  XNOR2X1 U1395 ( .A(n997), .B(n1), .Y(n979) );
  CLKAND2X4 U1396 ( .A(n167), .B(n254), .Y(n1236) );
  NOR2X1 U1397 ( .A(n226), .B(n169), .Y(n167) );
  XOR2X4 U1398 ( .A(n1232), .B(n72), .Y(product[27]) );
  XNOR2X4 U1399 ( .A(n203), .B(n74), .Y(product[25]) );
  CLKINVX4 U1400 ( .A(n224), .Y(n222) );
  NAND2X1 U1401 ( .A(n224), .B(n217), .Y(n215) );
  CLKINVX3 U1402 ( .A(n226), .Y(n224) );
  OAI22X1 U1403 ( .A0(n870), .A1(n40), .B0(n871), .B1(n41), .Y(n693) );
  OAI22X1 U1404 ( .A0(n1126), .A1(n41), .B0(n871), .B1(n40), .Y(n694) );
  OAI22X1 U1405 ( .A0(n915), .A1(n24), .B0(n914), .B1(n22), .Y(n736) );
  OAI22X1 U1406 ( .A0(n915), .A1(n22), .B0(n916), .B1(n24), .Y(n737) );
  OAI22X1 U1407 ( .A0(n1208), .A1(n53), .B0(n830), .B1(n51), .Y(n657) );
  ADDHX1 U1408 ( .A(n763), .B(n779), .CO(n600), .S(n601) );
  OAI22X1 U1409 ( .A0(n957), .A1(n9), .B0(n958), .B1(n11), .Y(n779) );
  OAI22X1 U1410 ( .A0(n894), .A1(n28), .B0(n895), .B1(n1016), .Y(n716) );
  AO21X1 U1411 ( .A0(n1016), .A1(n28), .B0(n894), .Y(n715) );
  XNOR2X1 U1412 ( .A(n984), .B(n25), .Y(n894) );
  BUFX12 U1413 ( .A(a[9]), .Y(n991) );
  OAI22X1 U1414 ( .A0(n962), .A1(n11), .B0(n961), .B1(n9), .Y(n783) );
  OAI22X1 U1415 ( .A0(n960), .A1(n9), .B0(n961), .B1(n11), .Y(n782) );
  ADDFHX2 U1416 ( .A(n630), .B(n767), .CI(n618), .CO(n615), .S(n616) );
  OAI22X1 U1417 ( .A0(n947), .A1(n15), .B0(n18), .B1(n1169), .Y(n630) );
  XNOR2X1 U1418 ( .A(n994), .B(n1), .Y(n976) );
  OAI22X1 U1419 ( .A0(n921), .A1(n1027), .B0(n1204), .B1(n23), .Y(n743) );
  ADDFHX2 U1420 ( .A(n747), .B(n628), .CI(n731), .CO(n598), .S(n599) );
  OAI22X1 U1421 ( .A0(n911), .A1(n28), .B0(n1016), .B1(n1036), .Y(n628) );
  OAI22X1 U1422 ( .A0(n929), .A1(n22), .B0(n24), .B1(n1196), .Y(n629) );
  XOR2X4 U1423 ( .A(n147), .B(n69), .Y(product[30]) );
  BUFX8 U1424 ( .A(a[11]), .Y(n989) );
  OAI22X1 U1425 ( .A0(n939), .A1(n15), .B0(n1207), .B1(n1018), .Y(n761) );
  XNOR2X1 U1426 ( .A(n995), .B(n25), .Y(n905) );
  XNOR2X4 U1427 ( .A(n232), .B(n77), .Y(product[22]) );
  XNOR2X1 U1428 ( .A(n995), .B(n19), .Y(n923) );
  XNOR2X1 U1429 ( .A(n994), .B(n7), .Y(n958) );
  OAI22X1 U1430 ( .A0(n971), .A1(n5), .B0(n970), .B1(n4), .Y(n792) );
  XNOR2X1 U1431 ( .A(n994), .B(n43), .Y(n850) );
  XNOR2X1 U1432 ( .A(n995), .B(n43), .Y(n851) );
  XNOR2X4 U1433 ( .A(n214), .B(n75), .Y(product[24]) );
  OAI22X1 U1434 ( .A0(n942), .A1(n1018), .B0(n941), .B1(n15), .Y(n763) );
  OAI22X1 U1435 ( .A0(n867), .A1(n40), .B0(n868), .B1(n41), .Y(n690) );
  OR2X1 U1436 ( .A(n948), .B(n9), .Y(n1210) );
  OR2XL U1437 ( .A(n949), .B(n12), .Y(n1211) );
  NAND2X1 U1438 ( .A(n1210), .B(n1211), .Y(n770) );
  OR2XL U1439 ( .A(n770), .B(n691), .Y(n517) );
  AO21X1 U1440 ( .A0(n18), .A1(n15), .B0(n930), .Y(n751) );
  XNOR2X1 U1441 ( .A(n984), .B(n13), .Y(n930) );
  OR2XL U1442 ( .A(n545), .B(n555), .Y(n1212) );
  CMPR42X2 U1443 ( .A(n561), .B(n551), .C(n558), .D(n548), .ICI(n554), .S(n545), .ICO(n543), .CO(n544) );
  CMPR42X2 U1444 ( .A(n566), .B(n562), .C(n567), .D(n563), .ICI(n559), .S(n556), .ICO(n554), .CO(n555) );
  NAND2XL U1445 ( .A(n986), .B(n25), .Y(n1214) );
  NAND2X1 U1446 ( .A(n1213), .B(n1036), .Y(n1215) );
  INVXL U1447 ( .A(n986), .Y(n1213) );
  BUFX12 U1448 ( .A(a[14]), .Y(n986) );
  OAI22X1 U1449 ( .A0(n895), .A1(n28), .B0(n896), .B1(n1016), .Y(n717) );
  BUFX12 U1450 ( .A(a[6]), .Y(n994) );
  XOR2X4 U1451 ( .A(n1228), .B(n76), .Y(product[23]) );
  OR2X2 U1452 ( .A(n886), .B(n1015), .Y(n1217) );
  NAND2X6 U1453 ( .A(n1216), .B(n1217), .Y(n707) );
  ADDFHX4 U1454 ( .A(n692), .B(n707), .CI(n677), .CO(n528), .S(n529) );
  XOR2X4 U1455 ( .A(n1237), .B(n73), .Y(product[26]) );
  NOR2BX2 U1456 ( .AN(n616), .B(n1219), .Y(n1218) );
  INVX8 U1457 ( .A(n166), .Y(n165) );
  AOI21X4 U1458 ( .A0(n110), .A1(n1137), .B0(n105), .Y(n103) );
  NAND2X2 U1459 ( .A(n109), .B(n1137), .Y(n102) );
  AO21XL U1460 ( .A0(n165), .A1(n123), .B0(n124), .Y(n1222) );
  CLKBUFX2 U1461 ( .A(n1021), .Y(n57) );
  OR2X1 U1462 ( .A(n884), .B(n34), .Y(n1221) );
  NAND2X2 U1463 ( .A(n1220), .B(n1221), .Y(n706) );
  ADDFHX2 U1464 ( .A(n676), .B(n706), .CI(n738), .CO(n515), .S(n516) );
  OR2X4 U1465 ( .A(n496), .B(n507), .Y(n1229) );
  OAI22XL U1466 ( .A0(n847), .A1(n48), .B0(n846), .B1(n46), .Y(n671) );
  NAND2X2 U1467 ( .A(n1226), .B(n1227), .Y(n448) );
  INVX1 U1468 ( .A(n448), .Y(n449) );
  XNOR2X1 U1469 ( .A(n787), .B(n771), .Y(n531) );
  NAND2XL U1470 ( .A(n990), .B(n43), .Y(n1224) );
  NAND2X1 U1471 ( .A(n1223), .B(n1033), .Y(n1225) );
  NAND2X1 U1472 ( .A(n1224), .B(n1225), .Y(n846) );
  INVXL U1473 ( .A(n990), .Y(n1223) );
  CMPR32X2 U1474 ( .A(n716), .B(n449), .C(n657), .CO(n446), .S(n447) );
  OR2X4 U1475 ( .A(n1230), .B(n1231), .Y(n771) );
  INVX1 U1476 ( .A(n468), .Y(n469) );
  CLKBUFX3 U1477 ( .A(n1017), .Y(n23) );
  OR2X2 U1478 ( .A(n815), .B(n59), .Y(n1226) );
  ADDFX2 U1479 ( .A(n699), .B(n448), .CI(n715), .CO(n438), .S(n439) );
  CLKINVX1 U1480 ( .A(n1229), .Y(n251) );
  INVX3 U1481 ( .A(n298), .Y(n296) );
  AO21X2 U1482 ( .A0(n1020), .A1(n4), .B0(n966), .Y(n787) );
  XNOR2X1 U1483 ( .A(n985), .B(n19), .Y(n913) );
  AOI21X2 U1484 ( .A0(n1136), .A1(n301), .B0(n296), .Y(n294) );
  OR2X1 U1485 ( .A(n787), .B(n771), .Y(n530) );
  NOR2BXL U1486 ( .AN(n61), .B(n57), .Y(n648) );
  CMPR42X2 U1487 ( .A(n753), .B(n769), .C(n675), .D(n690), .ICI(n647), .S(n505), .ICO(n503), .CO(n504) );
  XNOR2X1 U1488 ( .A(n998), .B(n7), .Y(n962) );
  INVXL U1489 ( .A(n49), .Y(n1032) );
  CLKXOR2X1 U1490 ( .A(b[4]), .B(b[5]), .Y(n1008) );
  XNOR2X1 U1491 ( .A(b[16]), .B(b[15]), .Y(n1022) );
  NOR2XL U1492 ( .A(n949), .B(n9), .Y(n1230) );
  CLKINVX4 U1493 ( .A(n283), .Y(n1241) );
  INVX4 U1494 ( .A(n292), .Y(n1244) );
  NOR2X4 U1495 ( .A(n145), .B(n138), .Y(n136) );
  NAND2X1 U1496 ( .A(n403), .B(n407), .Y(n146) );
  XNOR2X1 U1497 ( .A(n994), .B(n31), .Y(n886) );
  XOR2XL U1498 ( .A(b[14]), .B(b[15]), .Y(n1003) );
  NAND2XL U1499 ( .A(n985), .B(n13), .Y(n1234) );
  NAND2X1 U1500 ( .A(n1233), .B(n1169), .Y(n1235) );
  NAND2X1 U1501 ( .A(n1234), .B(n1235), .Y(n931) );
  INVXL U1502 ( .A(n985), .Y(n1233) );
  OAI22X1 U1503 ( .A0(n930), .A1(n15), .B0(n931), .B1(n18), .Y(n752) );
  OAI21X2 U1504 ( .A0(n315), .A1(n327), .B0(n316), .Y(n314) );
  AOI21X4 U1505 ( .A0(n162), .A1(n1127), .B0(n157), .Y(n155) );
  AOI21X4 U1506 ( .A0(n124), .A1(n1132), .B0(n119), .Y(n117) );
  OAI22X1 U1507 ( .A0(n888), .A1(n34), .B0(n1122), .B1(n1015), .Y(n710) );
  OAI22X1 U1508 ( .A0(n834), .A1(n51), .B0(n835), .B1(n53), .Y(n660) );
  NAND2X2 U1509 ( .A(n1238), .B(n1239), .Y(n492) );
  XNOR2XL U1510 ( .A(n990), .B(n25), .Y(n900) );
  XNOR2XL U1511 ( .A(n991), .B(n25), .Y(n901) );
  XNOR2XL U1512 ( .A(n998), .B(n37), .Y(n872) );
  XNOR2XL U1513 ( .A(n61), .B(n49), .Y(n838) );
  XNOR2XL U1514 ( .A(n988), .B(n25), .Y(n898) );
  XNOR2XL U1515 ( .A(n989), .B(n25), .Y(n899) );
  CLKBUFX2 U1516 ( .A(n1023), .Y(n46) );
  CLKBUFX4 U1517 ( .A(b[3]), .Y(n7) );
  XNOR2X2 U1518 ( .A(b[10]), .B(b[9]), .Y(n1025) );
  NOR2X6 U1519 ( .A(n1236), .B(n168), .Y(n166) );
  CMPR42X2 U1520 ( .A(n505), .B(n502), .C(n510), .D(n506), .ICI(n499), .S(n496), .ICO(n494), .CO(n495) );
  INVXL U1521 ( .A(n246), .Y(n240) );
  INVXL U1522 ( .A(n247), .Y(n241) );
  INVX1 U1523 ( .A(n272), .Y(n270) );
  BUFX2 U1524 ( .A(\product[39] ), .Y(\product[38] ) );
  NAND2XL U1525 ( .A(n370), .B(n249), .Y(n79) );
  INVXL U1526 ( .A(n248), .Y(n370) );
  INVXL U1527 ( .A(n289), .Y(n377) );
  INVXL U1528 ( .A(n311), .Y(n381) );
  XOR2X2 U1529 ( .A(n1240), .B(n85), .Y(product[14]) );
  CLKINVX1 U1530 ( .A(n107), .Y(n105) );
  OAI21X2 U1531 ( .A0(n333), .A1(n345), .B0(n334), .Y(n332) );
  NAND2X1 U1532 ( .A(n1134), .B(n331), .Y(n93) );
  NAND2X1 U1533 ( .A(n591), .B(n596), .Y(n309) );
  NAND2X1 U1534 ( .A(n556), .B(n564), .Y(n287) );
  NAND2X1 U1535 ( .A(n609), .B(n613), .Y(n325) );
  OAI22X2 U1536 ( .A0(n966), .A1(n4), .B0(n967), .B1(n1020), .Y(n788) );
  OAI22X2 U1537 ( .A0(n875), .A1(n40), .B0(n41), .B1(n1034), .Y(n626) );
  ADDFX2 U1538 ( .A(n711), .B(n626), .CI(n775), .CO(n569), .S(n570) );
  ADDFX2 U1539 ( .A(n744), .B(n728), .CI(n760), .CO(n579), .S(n580) );
  OAI22X1 U1540 ( .A0(n828), .A1(n53), .B0(n827), .B1(n51), .Y(n654) );
  OAI22XL U1541 ( .A0(n805), .A1(n58), .B0(n806), .B1(n1011), .Y(n634) );
  XNOR2X1 U1542 ( .A(n997), .B(n49), .Y(n835) );
  XNOR2X1 U1543 ( .A(n997), .B(n43), .Y(n853) );
  XNOR2X1 U1544 ( .A(n988), .B(n19), .Y(n916) );
  XNOR2X1 U1545 ( .A(n989), .B(n19), .Y(n917) );
  XNOR2X1 U1546 ( .A(n985), .B(n1), .Y(n967) );
  XNOR2XL U1547 ( .A(n992), .B(n1), .Y(n974) );
  NAND2BXL U1548 ( .AN(n61), .B(n25), .Y(n911) );
  XNOR2XL U1549 ( .A(n990), .B(n49), .Y(n828) );
  BUFX8 U1550 ( .A(a[4]), .Y(n996) );
  NAND2X2 U1551 ( .A(n1003), .B(n1023), .Y(n1013) );
  XNOR2X2 U1552 ( .A(b[12]), .B(b[11]), .Y(n1024) );
  OR2X2 U1553 ( .A(n851), .B(n47), .Y(n1238) );
  OR2X2 U1554 ( .A(n850), .B(n46), .Y(n1239) );
  INVXL U1555 ( .A(n220), .Y(n218) );
  INVXL U1556 ( .A(n238), .Y(n236) );
  NOR2XL U1557 ( .A(n150), .B(n143), .Y(n141) );
  INVXL U1558 ( .A(n237), .Y(n235) );
  AO21X4 U1559 ( .A0(n1241), .A1(n1242), .B0(n1243), .Y(n254) );
  AOI21X2 U1560 ( .A0(n1135), .A1(n323), .B0(n318), .Y(n316) );
  NAND2X2 U1561 ( .A(n1135), .B(n1128), .Y(n315) );
  OA21X4 U1562 ( .A0(n1244), .A1(n1245), .B0(n1246), .Y(n283) );
  INVX3 U1563 ( .A(n191), .Y(n189) );
  NAND2XL U1564 ( .A(n377), .B(n290), .Y(n86) );
  NAND2XL U1565 ( .A(n381), .B(n312), .Y(n90) );
  INVX3 U1566 ( .A(n159), .Y(n157) );
  INVXL U1567 ( .A(n281), .Y(n279) );
  OAI21X4 U1568 ( .A0(n305), .A1(n293), .B0(n294), .Y(n292) );
  AOI21X2 U1569 ( .A0(n350), .A1(n1133), .B0(n347), .Y(n345) );
  AOI21X2 U1570 ( .A0(n332), .A1(n1134), .B0(n329), .Y(n327) );
  CMPR42X2 U1571 ( .A(n488), .B(n478), .C(n475), .D(n485), .ICI(n481), .S(n472), .ICO(n470), .CO(n471) );
  NOR2X1 U1572 ( .A(n545), .B(n555), .Y(n280) );
  ADDHX1 U1573 ( .A(n799), .B(n783), .CO(n617), .S(n618) );
  CMPR42X2 U1574 ( .A(n668), .B(n640), .C(n428), .D(n423), .ICI(n424), .S(n420), .ICO(n418), .CO(n419) );
  CMPR42X2 U1575 ( .A(n683), .B(n655), .C(n429), .D(n436), .ICI(n432), .S(n426), .ICO(n424), .CO(n425) );
  CMPR42X2 U1576 ( .A(n480), .B(n490), .C(n487), .D(n719), .ICI(n484), .S(n475), .ICO(n473), .CO(n474) );
  CMPR42X2 U1577 ( .A(n431), .B(n641), .C(n669), .D(n438), .ICI(n435), .S(n429), .ICO(n427), .CO(n428) );
  INVX3 U1578 ( .A(n430), .Y(n431) );
  CMPR42X2 U1579 ( .A(n514), .B(n526), .C(n523), .D(n511), .ICI(n519), .S(n508), .ICO(n506), .CO(n507) );
  AO21XL U1580 ( .A0(n24), .A1(n22), .B0(n912), .Y(n733) );
  ADDHX1 U1581 ( .A(n789), .B(n709), .CO(n552), .S(n553) );
  AO21XL U1582 ( .A0(n41), .A1(n40), .B0(n858), .Y(n681) );
  ADDFX1 U1583 ( .A(n417), .B(n653), .CI(n421), .CO(n414), .S(n415) );
  OAI22X1 U1584 ( .A0(n954), .A1(n12), .B0(n953), .B1(n1029), .Y(n775) );
  CMPR42X2 U1585 ( .A(n739), .B(n663), .C(n529), .D(n755), .ICI(n723), .S(n524), .ICO(n522), .CO(n523) );
  AO21XL U1586 ( .A0(n36), .A1(n34), .B0(n1123), .Y(n698) );
  AO21XL U1587 ( .A0(n12), .A1(n9), .B0(n948), .Y(n769) );
  NAND2BXL U1588 ( .AN(n353), .B(n354), .Y(n98) );
  ADDFXL U1589 ( .A(n634), .B(n396), .CI(n649), .CO(n392), .S(n393) );
  AO21XL U1590 ( .A0(n53), .A1(n51), .B0(n822), .Y(n649) );
  OAI22X1 U1591 ( .A0(n804), .A1(n58), .B0(n805), .B1(n1011), .Y(n390) );
  AO21XL U1592 ( .A0(n1011), .A1(n58), .B0(n804), .Y(n633) );
  NAND2BXL U1593 ( .AN(n61), .B(n7), .Y(n965) );
  XNOR2XL U1594 ( .A(n985), .B(n31), .Y(n877) );
  XNOR2XL U1595 ( .A(n984), .B(n31), .Y(n876) );
  XNOR2XL U1596 ( .A(n999), .B(n25), .Y(n909) );
  XNOR2XL U1597 ( .A(n999), .B(n31), .Y(n891) );
  XNOR2XL U1598 ( .A(n999), .B(n43), .Y(n855) );
  XNOR2XL U1599 ( .A(n985), .B(n25), .Y(n895) );
  XNOR2XL U1600 ( .A(n990), .B(n37), .Y(n864) );
  XNOR2XL U1601 ( .A(n989), .B(n43), .Y(n845) );
  XNOR2XL U1602 ( .A(n989), .B(n37), .Y(n863) );
  XNOR2XL U1603 ( .A(n990), .B(n31), .Y(n882) );
  XNOR2XL U1604 ( .A(n998), .B(n25), .Y(n908) );
  XNOR2XL U1605 ( .A(n993), .B(n49), .Y(n831) );
  XNOR2XL U1606 ( .A(n993), .B(n37), .Y(n867) );
  XNOR2XL U1607 ( .A(n998), .B(n55), .Y(n818) );
  XNOR2XL U1608 ( .A(n993), .B(n43), .Y(n849) );
  XNOR2XL U1609 ( .A(n984), .B(n37), .Y(n858) );
  XNOR2XL U1610 ( .A(n984), .B(n19), .Y(n912) );
  XNOR2XL U1611 ( .A(n61), .B(n25), .Y(n910) );
  XNOR2XL U1612 ( .A(n61), .B(n19), .Y(n928) );
  XNOR2XL U1613 ( .A(n61), .B(n43), .Y(n856) );
  XNOR2XL U1614 ( .A(n61), .B(n55), .Y(n820) );
  NAND2BXL U1615 ( .AN(n61), .B(n13), .Y(n947) );
  NAND2BXL U1616 ( .AN(n61), .B(n37), .Y(n875) );
  NAND2BXL U1617 ( .AN(n61), .B(n19), .Y(n929) );
  NAND2BXL U1618 ( .AN(n61), .B(n31), .Y(n893) );
  NAND2BXL U1619 ( .AN(n61), .B(n49), .Y(n839) );
  NAND2BXL U1620 ( .AN(n61), .B(n43), .Y(n857) );
  XNOR2XL U1621 ( .A(n984), .B(n43), .Y(n840) );
  XNOR2XL U1622 ( .A(n988), .B(n37), .Y(n862) );
  XNOR2XL U1623 ( .A(n992), .B(n55), .Y(n812) );
  XNOR2XL U1624 ( .A(n992), .B(n13), .Y(n938) );
  XNOR2XL U1625 ( .A(n999), .B(n55), .Y(n819) );
  XNOR2XL U1626 ( .A(n997), .B(n55), .Y(n817) );
  XNOR2XL U1627 ( .A(n992), .B(n49), .Y(n830) );
  XNOR2XL U1628 ( .A(n992), .B(n25), .Y(n902) );
  XNOR2XL U1629 ( .A(n988), .B(n31), .Y(n880) );
  XNOR2XL U1630 ( .A(n992), .B(n19), .Y(n920) );
  XNOR2XL U1631 ( .A(n992), .B(n37), .Y(n866) );
  XNOR2XL U1632 ( .A(n992), .B(n43), .Y(n848) );
  XNOR2XL U1633 ( .A(n990), .B(n55), .Y(n810) );
  XNOR2XL U1634 ( .A(n989), .B(n55), .Y(n809) );
  XNOR2XL U1635 ( .A(n989), .B(n49), .Y(n827) );
  XNOR2XL U1636 ( .A(n989), .B(n31), .Y(n881) );
  XNOR2XL U1637 ( .A(n987), .B(n37), .Y(n861) );
  XNOR2XL U1638 ( .A(n987), .B(n25), .Y(n897) );
  XNOR2XL U1639 ( .A(n991), .B(n13), .Y(n937) );
  XNOR2XL U1640 ( .A(n991), .B(n49), .Y(n829) );
  XNOR2XL U1641 ( .A(n991), .B(n19), .Y(n919) );
  XNOR2XL U1642 ( .A(n991), .B(n31), .Y(n883) );
  XNOR2XL U1643 ( .A(n991), .B(n37), .Y(n865) );
  XNOR2XL U1644 ( .A(n986), .B(n55), .Y(n806) );
  XNOR2XL U1645 ( .A(n988), .B(n55), .Y(n808) );
  XNOR2XL U1646 ( .A(n986), .B(n49), .Y(n824) );
  XNOR2XL U1647 ( .A(n985), .B(n49), .Y(n823) );
  XNOR2XL U1648 ( .A(n987), .B(n55), .Y(n807) );
  XNOR2XL U1649 ( .A(n991), .B(n55), .Y(n811) );
  XNOR2XL U1650 ( .A(n987), .B(n49), .Y(n825) );
  XNOR2XL U1651 ( .A(n991), .B(n43), .Y(n847) );
  XNOR2XL U1652 ( .A(n984), .B(n49), .Y(n822) );
  CLKBUFX2 U1653 ( .A(n1021), .Y(n58) );
  XNOR2X1 U1654 ( .A(b[8]), .B(b[7]), .Y(n1026) );
  XNOR2X1 U1655 ( .A(b[4]), .B(b[3]), .Y(n1028) );
  NAND2X4 U1656 ( .A(n1009), .B(n1029), .Y(n1019) );
  INVX1 U1657 ( .A(b[0]), .Y(n1030) );
  CLKINVX1 U1658 ( .A(n211), .Y(n209) );
  CLKINVX1 U1659 ( .A(n152), .Y(n150) );
  NOR2X1 U1660 ( .A(n150), .B(n134), .Y(n132) );
  NAND2X1 U1661 ( .A(n246), .B(n235), .Y(n233) );
  CLKINVX1 U1662 ( .A(n116), .Y(n114) );
  NAND2X1 U1663 ( .A(n366), .B(n213), .Y(n75) );
  CLKINVX1 U1664 ( .A(n212), .Y(n366) );
  NAND2X1 U1665 ( .A(n368), .B(n231), .Y(n77) );
  CLKINVX1 U1666 ( .A(n230), .Y(n368) );
  AOI21X1 U1667 ( .A0(n225), .A1(n217), .B0(n218), .Y(n216) );
  AOI21X1 U1668 ( .A0(n247), .A1(n235), .B0(n236), .Y(n234) );
  AOI21X1 U1669 ( .A0(n225), .A1(n182), .B0(n183), .Y(n181) );
  NAND2X1 U1670 ( .A(n374), .B(n276), .Y(n83) );
  AOI21X1 U1671 ( .A0(n1125), .A1(n1212), .B0(n279), .Y(n277) );
  CLKINVX1 U1672 ( .A(n275), .Y(n374) );
  CLKINVX1 U1673 ( .A(n273), .Y(n271) );
  CLKINVX1 U1674 ( .A(n274), .Y(n272) );
  NOR2X1 U1675 ( .A(n271), .B(n264), .Y(n262) );
  CLKINVX1 U1676 ( .A(n137), .Y(n135) );
  CLKINVX1 U1677 ( .A(n136), .Y(n134) );
  CLKINVX1 U1678 ( .A(n365), .Y(n197) );
  CLKINVX1 U1679 ( .A(n117), .Y(n115) );
  XNOR2X1 U1680 ( .A(n326), .B(n92), .Y(product[7]) );
  NAND2X1 U1681 ( .A(n1128), .B(n325), .Y(n92) );
  NAND2X1 U1682 ( .A(n1129), .B(n164), .Y(n71) );
  NAND2X1 U1683 ( .A(n1130), .B(n178), .Y(n72) );
  NAND2X1 U1684 ( .A(n364), .B(n191), .Y(n73) );
  CLKINVX1 U1685 ( .A(n190), .Y(n364) );
  NAND2X1 U1686 ( .A(n376), .B(n287), .Y(n85) );
  CLKINVX1 U1687 ( .A(n286), .Y(n376) );
  NAND2X1 U1688 ( .A(n380), .B(n309), .Y(n89) );
  CLKINVX1 U1689 ( .A(n308), .Y(n380) );
  XNOR2X1 U1690 ( .A(n1125), .B(n84), .Y(product[15]) );
  NAND2X1 U1691 ( .A(n1212), .B(n281), .Y(n84) );
  NOR2X1 U1692 ( .A(n308), .B(n311), .Y(n306) );
  NOR2X2 U1693 ( .A(n534), .B(n544), .Y(n275) );
  CLKINVX1 U1694 ( .A(n130), .Y(n128) );
  NAND2X1 U1695 ( .A(n1137), .B(n107), .Y(n64) );
  CLKINVX1 U1696 ( .A(n178), .Y(n176) );
  XOR2X1 U1697 ( .A(n321), .B(n91), .Y(product[8]) );
  NAND2X1 U1698 ( .A(n1135), .B(n320), .Y(n91) );
  AOI21X1 U1699 ( .A0(n326), .A1(n1128), .B0(n323), .Y(n321) );
  XOR2X1 U1700 ( .A(n291), .B(n86), .Y(product[13]) );
  NAND2X1 U1701 ( .A(n372), .B(n260), .Y(n81) );
  CLKINVX1 U1702 ( .A(n259), .Y(n372) );
  NAND2X1 U1703 ( .A(n265), .B(n267), .Y(n82) );
  AOI21X1 U1704 ( .A0(n1125), .A1(n273), .B0(n270), .Y(n268) );
  XOR2X1 U1705 ( .A(n313), .B(n90), .Y(product[9]) );
  NAND2X1 U1706 ( .A(n356), .B(n112), .Y(n65) );
  AOI21X1 U1707 ( .A0(n165), .A1(n114), .B0(n115), .Y(n113) );
  CLKINVX1 U1708 ( .A(n111), .Y(n356) );
  NAND2X1 U1709 ( .A(n1131), .B(n130), .Y(n67) );
  NAND2X1 U1710 ( .A(n359), .B(n139), .Y(n68) );
  AOI21X1 U1711 ( .A0(n165), .A1(n141), .B0(n142), .Y(n140) );
  CLKINVX1 U1712 ( .A(n138), .Y(n359) );
  NAND2X1 U1713 ( .A(n1127), .B(n159), .Y(n70) );
  AOI21X1 U1714 ( .A0(n165), .A1(n1129), .B0(n162), .Y(n160) );
  NAND2X1 U1715 ( .A(n144), .B(n146), .Y(n69) );
  AOI21X1 U1716 ( .A0(n165), .A1(n152), .B0(n153), .Y(n147) );
  XOR2X1 U1717 ( .A(n253), .B(n80), .Y(product[19]) );
  NAND2X1 U1718 ( .A(n1229), .B(n252), .Y(n80) );
  NAND2X1 U1719 ( .A(n461), .B(n471), .Y(n231) );
  NAND2X1 U1720 ( .A(n534), .B(n544), .Y(n276) );
  CLKINVX1 U1721 ( .A(n292), .Y(n291) );
  CLKINVX1 U1722 ( .A(n265), .Y(n264) );
  CLKINVX1 U1723 ( .A(n266), .Y(n265) );
  CLKINVX1 U1724 ( .A(n327), .Y(n326) );
  CLKINVX1 U1725 ( .A(n325), .Y(n323) );
  CLKINVX1 U1726 ( .A(n164), .Y(n162) );
  OAI21XL U1727 ( .A0(n155), .A1(n143), .B0(n146), .Y(n142) );
  CLKINVX1 U1728 ( .A(n144), .Y(n143) );
  CLKINVX1 U1729 ( .A(n145), .Y(n144) );
  CLKINVX1 U1730 ( .A(n345), .Y(n344) );
  XNOR2X1 U1731 ( .A(n332), .B(n93), .Y(product[6]) );
  XNOR2X1 U1732 ( .A(n304), .B(n88), .Y(product[11]) );
  NAND2X1 U1733 ( .A(n300), .B(n303), .Y(n88) );
  NAND2X1 U1734 ( .A(n1136), .B(n300), .Y(n293) );
  CLKINVX1 U1735 ( .A(n349), .Y(n347) );
  NOR2X2 U1736 ( .A(n556), .B(n564), .Y(n286) );
  NOR2X2 U1737 ( .A(n591), .B(n596), .Y(n308) );
  AOI21X1 U1738 ( .A0(n335), .A1(n341), .B0(n1218), .Y(n334) );
  NAND2X1 U1739 ( .A(n335), .B(n386), .Y(n333) );
  NAND2X1 U1740 ( .A(n545), .B(n555), .Y(n281) );
  NAND2X1 U1741 ( .A(n1136), .B(n298), .Y(n87) );
  AOI21X1 U1742 ( .A0(n304), .A1(n300), .B0(n301), .Y(n299) );
  NAND2X1 U1743 ( .A(n565), .B(n574), .Y(n290) );
  NAND2X1 U1744 ( .A(n802), .B(n786), .Y(n352) );
  NAND2X1 U1745 ( .A(n604), .B(n608), .Y(n320) );
  NAND2X1 U1746 ( .A(n420), .B(n425), .Y(n178) );
  NAND2X1 U1747 ( .A(n412), .B(n408), .Y(n159) );
  NAND2X1 U1748 ( .A(n433), .B(n426), .Y(n191) );
  NAND2X1 U1749 ( .A(n508), .B(n520), .Y(n260) );
  XNOR2X1 U1750 ( .A(n96), .B(n350), .Y(product[3]) );
  NAND2X1 U1751 ( .A(n1133), .B(n349), .Y(n96) );
  NAND2X1 U1752 ( .A(n386), .B(n343), .Y(n95) );
  CLKINVX1 U1753 ( .A(n342), .Y(n386) );
  XOR2X1 U1754 ( .A(n97), .B(n354), .Y(product[2]) );
  NAND2X1 U1755 ( .A(n388), .B(n352), .Y(n97) );
  CLKINVX1 U1756 ( .A(n351), .Y(n388) );
  NAND2X1 U1757 ( .A(n335), .B(n338), .Y(n94) );
  AOI21X1 U1758 ( .A0(n344), .A1(n386), .B0(n341), .Y(n339) );
  NAND2X1 U1759 ( .A(n399), .B(n395), .Y(n130) );
  NAND2X1 U1760 ( .A(n400), .B(n402), .Y(n139) );
  NAND2X1 U1761 ( .A(n633), .B(n390), .Y(n107) );
  NAND2X1 U1762 ( .A(n394), .B(n393), .Y(n121) );
  CLKINVX1 U1763 ( .A(n390), .Y(n391) );
  NAND2X1 U1764 ( .A(n392), .B(n391), .Y(n112) );
  OAI22X1 U1765 ( .A0(n1123), .A1(n34), .B0(n1209), .B1(n36), .Y(n430) );
  CMPR42X1 U1766 ( .A(n798), .B(n782), .C(n750), .D(n766), .ICI(n617), .S(n614), .ICO(n612), .CO(n613) );
  NOR2BX1 U1767 ( .AN(n61), .B(n1027), .Y(n750) );
  OAI22XL U1768 ( .A0(n944), .A1(n15), .B0(n945), .B1(n1018), .Y(n766) );
  CMPR42X1 U1769 ( .A(n580), .B(n584), .C(n578), .D(n585), .ICI(n581), .S(n575), .ICO(n573), .CO(n574) );
  CMPR42X1 U1770 ( .A(n730), .B(n598), .C(n794), .D(n595), .ICI(n594), .S(n591), .ICO(n589), .CO(n590) );
  OAI22XL U1771 ( .A0(n908), .A1(n28), .B0(n909), .B1(n29), .Y(n730) );
  OAI22XL U1772 ( .A0(n937), .A1(n15), .B0(n938), .B1(n1018), .Y(n759) );
  OAI22XL U1773 ( .A0(n969), .A1(n4), .B0(n970), .B1(n5), .Y(n791) );
  OAI22XL U1774 ( .A0(n811), .A1(n58), .B0(n812), .B1(n59), .Y(n640) );
  OAI22XL U1775 ( .A0(n861), .A1(n40), .B0(n862), .B1(n41), .Y(n684) );
  OAI22XL U1776 ( .A0(n810), .A1(n59), .B0(n809), .B1(n58), .Y(n638) );
  OAI22XL U1777 ( .A0(n825), .A1(n51), .B0(n826), .B1(n53), .Y(n652) );
  OAI22XL U1778 ( .A0(n811), .A1(n59), .B0(n810), .B1(n58), .Y(n639) );
  OAI22XL U1779 ( .A0(n829), .A1(n53), .B0(n828), .B1(n51), .Y(n655) );
  OAI22XL U1780 ( .A0(n836), .A1(n53), .B0(n835), .B1(n51), .Y(n661) );
  OAI22XL U1781 ( .A0(n912), .A1(n22), .B0(n913), .B1(n24), .Y(n734) );
  OAI22XL U1782 ( .A0(n818), .A1(n57), .B0(n819), .B1(n59), .Y(n646) );
  NOR2X2 U1783 ( .A(n583), .B(n590), .Y(n302) );
  NOR2X2 U1784 ( .A(n616), .B(n619), .Y(n337) );
  OAI22XL U1785 ( .A0(n882), .A1(n36), .B0(n881), .B1(n34), .Y(n703) );
  CMPR42X1 U1786 ( .A(n682), .B(n430), .C(n698), .D(n654), .ICI(n427), .S(n423), .ICO(n421), .CO(n422) );
  NOR2BX1 U1787 ( .AN(n61), .B(n15), .Y(n768) );
  OAI22XL U1788 ( .A0(n962), .A1(n9), .B0(n963), .B1(n11), .Y(n784) );
  OAI22XL U1789 ( .A0(n849), .A1(n1023), .B0(n850), .B1(n47), .Y(n674) );
  OAI22XL U1790 ( .A0(n865), .A1(n40), .B0(n866), .B1(n41), .Y(n688) );
  OAI22XL U1791 ( .A0(n818), .A1(n59), .B0(n817), .B1(n57), .Y(n645) );
  CMPR42X1 U1792 ( .A(n648), .B(n662), .C(n530), .D(n518), .ICI(n525), .S(n514), .ICO(n512), .CO(n513) );
  XNOR2X1 U1793 ( .A(n770), .B(n691), .Y(n518) );
  CMPR42X1 U1794 ( .A(n734), .B(n469), .C(n673), .D(n702), .ICI(n476), .S(n467), .ICO(n465), .CO(n466) );
  OAI22XL U1795 ( .A0(n881), .A1(n36), .B0(n880), .B1(n34), .Y(n702) );
  CMPR42X1 U1796 ( .A(n517), .B(n661), .C(n623), .D(n721), .ICI(n705), .S(n502), .ICO(n500), .CO(n501) );
  OAI22XL U1797 ( .A0(n883), .A1(n34), .B0(n884), .B1(n1015), .Y(n705) );
  OAI22XL U1798 ( .A0(n900), .A1(n1016), .B0(n899), .B1(n28), .Y(n721) );
  NAND2X1 U1799 ( .A(n614), .B(n615), .Y(n331) );
  NAND2X1 U1800 ( .A(n583), .B(n590), .Y(n303) );
  NAND2X1 U1801 ( .A(n575), .B(n582), .Y(n298) );
  CMPR42X1 U1802 ( .A(n697), .B(n792), .C(n712), .D(n587), .ICI(n776), .S(n578), .ICO(n576), .CO(n577) );
  NOR2BX1 U1803 ( .AN(n61), .B(n40), .Y(n697) );
  OAI22XL U1804 ( .A0(n813), .A1(n59), .B0(n812), .B1(n57), .Y(n641) );
  CMPR42X1 U1805 ( .A(n642), .B(n670), .C(n439), .D(n446), .ICI(n656), .S(n437), .ICO(n435), .CO(n436) );
  OAI22XL U1806 ( .A0(n813), .A1(n57), .B0(n814), .B1(n59), .Y(n642) );
  OAI22XL U1807 ( .A0(n829), .A1(n51), .B0(n830), .B1(n53), .Y(n656) );
  CMPR42X1 U1808 ( .A(n732), .B(n748), .C(n610), .D(n606), .ICI(n607), .S(n604), .ICO(n602), .CO(n603) );
  NOR2BX1 U1809 ( .AN(n61), .B(n28), .Y(n732) );
  OAI22XL U1810 ( .A0(n883), .A1(n36), .B0(n882), .B1(n34), .Y(n704) );
  OAI22XL U1811 ( .A0(n919), .A1(n22), .B0(n920), .B1(n23), .Y(n741) );
  OAI22XL U1812 ( .A0(n856), .A1(n47), .B0(n855), .B1(n1023), .Y(n679) );
  OAI22XL U1813 ( .A0(n953), .A1(n12), .B0(n952), .B1(n9), .Y(n774) );
  OAI22XL U1814 ( .A0(n901), .A1(n28), .B0(n902), .B1(n29), .Y(n723) );
  CMPR42X1 U1815 ( .A(n515), .B(n512), .C(n737), .D(n509), .ICI(n513), .S(n499), .ICO(n497), .CO(n498) );
  OAI22XL U1816 ( .A0(n937), .A1(n18), .B0(n936), .B1(n15), .Y(n758) );
  NOR2BX1 U1817 ( .AN(n61), .B(n1023), .Y(n680) );
  NOR2BX1 U1818 ( .AN(n61), .B(n34), .Y(n714) );
  CMPR42X1 U1819 ( .A(n625), .B(n757), .C(n560), .D(n773), .ICI(n557), .S(n548), .ICO(n546), .CO(n547) );
  OAI22XL U1820 ( .A0(n857), .A1(n46), .B0(n48), .B1(n1033), .Y(n625) );
  CMPR42X1 U1821 ( .A(n685), .B(n456), .C(n447), .D(n700), .ICI(n671), .S(n445), .ICO(n443), .CO(n444) );
  OAI22XL U1822 ( .A0(n863), .A1(n41), .B0(n862), .B1(n40), .Y(n685) );
  OAI22XL U1823 ( .A0(n847), .A1(n46), .B0(n848), .B1(n47), .Y(n672) );
  OAI22XL U1824 ( .A0(n816), .A1(n57), .B0(n817), .B1(n59), .Y(n644) );
  OAI22XL U1825 ( .A0(n865), .A1(n41), .B0(n864), .B1(n40), .Y(n687) );
  NAND2X1 U1826 ( .A(n620), .B(n621), .Y(n343) );
  OAI22XL U1827 ( .A0(n919), .A1(n24), .B0(n918), .B1(n22), .Y(n740) );
  OAI22XL U1828 ( .A0(n901), .A1(n1016), .B0(n900), .B1(n28), .Y(n722) );
  CMPR42X1 U1829 ( .A(n601), .B(n605), .C(n602), .D(n795), .ICI(n599), .S(n597), .ICO(n595), .CO(n596) );
  OAI22XL U1830 ( .A0(n973), .A1(n4), .B0(n974), .B1(n5), .Y(n795) );
  OAI22XL U1831 ( .A0(n820), .A1(n59), .B0(n819), .B1(n57), .Y(n647) );
  OAI22XL U1832 ( .A0(n816), .A1(n59), .B0(n815), .B1(n57), .Y(n643) );
  CMPR42X1 U1833 ( .A(n664), .B(n542), .C(n549), .D(n772), .ICI(n546), .S(n537), .ICO(n535), .CO(n536) );
  NOR2BX1 U1834 ( .AN(n61), .B(n51), .Y(n664) );
  OAI22XL U1835 ( .A0(n939), .A1(n1018), .B0(n938), .B1(n15), .Y(n760) );
  OAI22XL U1836 ( .A0(n822), .A1(n51), .B0(n823), .B1(n53), .Y(n396) );
  OAI22X1 U1837 ( .A0(n840), .A1(n46), .B0(n841), .B1(n48), .Y(n404) );
  NOR2BX1 U1838 ( .AN(n61), .B(n1030), .Y(product[0]) );
  AO21X1 U1839 ( .A0(n48), .A1(n46), .B0(n840), .Y(n665) );
  OAI22XL U1840 ( .A0(n823), .A1(n51), .B0(n1121), .B1(n53), .Y(n650) );
  OAI22XL U1841 ( .A0(n807), .A1(n58), .B0(n808), .B1(n59), .Y(n636) );
  OAI22XL U1842 ( .A0(n809), .A1(n59), .B0(n808), .B1(n58), .Y(n637) );
  CLKINVX1 U1843 ( .A(n404), .Y(n405) );
  OAI22XL U1844 ( .A0(n825), .A1(n53), .B0(n1121), .B1(n51), .Y(n651) );
  ADDFX2 U1845 ( .A(n397), .B(n398), .CI(n635), .CO(n394), .S(n395) );
  CLKINVX1 U1846 ( .A(n396), .Y(n397) );
  OAI22XL U1847 ( .A0(n807), .A1(n1011), .B0(n806), .B1(n58), .Y(n635) );
  CLKINVX1 U1848 ( .A(n98), .Y(product[1]) );
  XNOR2X1 U1849 ( .A(n61), .B(n1), .Y(n982) );
  XNOR2X1 U1850 ( .A(n61), .B(n7), .Y(n964) );
  CMPR42X1 U1851 ( .A(n793), .B(n713), .C(n593), .D(n589), .ICI(n586), .S(n583), .ICO(n581), .CO(n582) );
  OAI22XL U1852 ( .A0(n892), .A1(n1015), .B0(n891), .B1(n1025), .Y(n713) );
  XNOR2X1 U1853 ( .A(n61), .B(n31), .Y(n892) );
  XNOR2X1 U1854 ( .A(n996), .B(n13), .Y(n942) );
  XNOR2X1 U1855 ( .A(n993), .B(n1), .Y(n975) );
  XNOR2X1 U1856 ( .A(n996), .B(n7), .Y(n960) );
  XNOR2X1 U1857 ( .A(n996), .B(n49), .Y(n834) );
  XNOR2X1 U1858 ( .A(n996), .B(n43), .Y(n852) );
  XNOR2X1 U1859 ( .A(n996), .B(n31), .Y(n888) );
  XNOR2X1 U1860 ( .A(n996), .B(n19), .Y(n924) );
  XNOR2X1 U1861 ( .A(n996), .B(n37), .Y(n870) );
  XNOR2X1 U1862 ( .A(n996), .B(n25), .Y(n906) );
  XNOR2X1 U1863 ( .A(n987), .B(n31), .Y(n879) );
  XNOR2X1 U1864 ( .A(n996), .B(n55), .Y(n816) );
  XNOR2X1 U1865 ( .A(n993), .B(n7), .Y(n957) );
  XNOR2X1 U1866 ( .A(n996), .B(n1), .Y(n978) );
  XNOR2X1 U1867 ( .A(n995), .B(n1), .Y(n977) );
  XNOR2X1 U1868 ( .A(n989), .B(n7), .Y(n953) );
  XNOR2X1 U1869 ( .A(n999), .B(n1), .Y(n981) );
  XNOR2X1 U1870 ( .A(n999), .B(n13), .Y(n945) );
  XNOR2X1 U1871 ( .A(n997), .B(n13), .Y(n943) );
  XNOR2X1 U1872 ( .A(n992), .B(n31), .Y(n884) );
  XNOR2X1 U1873 ( .A(n999), .B(n7), .Y(n963) );
  XNOR2X1 U1874 ( .A(n984), .B(n1), .Y(n966) );
  OAI22XL U1875 ( .A0(n821), .A1(n58), .B0(n59), .B1(n1146), .Y(n623) );
  NAND2BX1 U1876 ( .AN(n61), .B(n55), .Y(n821) );
  XNOR2X1 U1877 ( .A(n61), .B(n37), .Y(n874) );
  XNOR2X1 U1878 ( .A(n985), .B(n55), .Y(n805) );
  XNOR2X1 U1879 ( .A(n984), .B(n55), .Y(n804) );
  CLKBUFX3 U1880 ( .A(n1027), .Y(n22) );
  CLKBUFX3 U1881 ( .A(n1025), .Y(n34) );
  CLKBUFX3 U1882 ( .A(n1026), .Y(n28) );
  CLKBUFX3 U1883 ( .A(n1024), .Y(n40) );
  CLKBUFX3 U1884 ( .A(n1030), .Y(n4) );
  CLKBUFX3 U1885 ( .A(n1022), .Y(n51) );
  CLKBUFX3 U1886 ( .A(n1029), .Y(n9) );
  CLKBUFX3 U1887 ( .A(n1028), .Y(n15) );
  CLKBUFX3 U1888 ( .A(n1016), .Y(n29) );
  CLKBUFX3 U1889 ( .A(n1019), .Y(n11) );
  CLKBUFX3 U1890 ( .A(n1018), .Y(n18) );
  CLKBUFX3 U1891 ( .A(n1017), .Y(n24) );
  CLKBUFX3 U1892 ( .A(n1015), .Y(n36) );
  CLKBUFX3 U1893 ( .A(n1013), .Y(n48) );
  CLKINVX1 U1894 ( .A(n37), .Y(n1034) );
  CLKINVX1 U1895 ( .A(n43), .Y(n1033) );
  CLKINVX1 U1896 ( .A(n25), .Y(n1036) );
  XNOR2X2 U1897 ( .A(b[18]), .B(b[17]), .Y(n1021) );
  XNOR2X2 U1898 ( .A(b[14]), .B(b[13]), .Y(n1023) );
  XOR2X1 U1899 ( .A(b[18]), .B(b[19]), .Y(n1001) );
  NAND2X1 U1900 ( .A(n1004), .B(n1024), .Y(n1014) );
  XOR2X1 U1901 ( .A(b[12]), .B(b[13]), .Y(n1004) );
  NAND2X1 U1902 ( .A(n1002), .B(n1022), .Y(n1012) );
  XOR2X1 U1903 ( .A(b[16]), .B(b[17]), .Y(n1002) );
  XOR2X1 U1904 ( .A(b[2]), .B(b[3]), .Y(n1009) );
  NAND2X1 U1905 ( .A(n1007), .B(n1027), .Y(n1017) );
  XOR2X1 U1906 ( .A(b[6]), .B(b[7]), .Y(n1007) );
  XOR2X1 U1907 ( .A(b[8]), .B(b[9]), .Y(n1006) );
  NAND2X1 U1908 ( .A(n1010), .B(n1030), .Y(n1020) );
  XOR2X1 U1909 ( .A(b[0]), .B(b[1]), .Y(n1010) );
endmodule


module CONV_DW01_add_5 ( A, B, CI, SUM, CO );
  input [43:0] A;
  input [43:0] B;
  output [43:0] SUM;
  input CI;
  output CO;
  wire   n2, n3, n4, n5, n6, n7, n8, n9, n10, n11, n12, n13, n14, n15, n16,
         n17, n18, n19, n20, n21, n22, n23, n24, n25, n26, n27, n28, n29, n30,
         n31, n32, n33, n34, n35, n36, n37, n38, n39, n40, n41, n42, n43, n44,
         n45, n47, n48, n53, n54, n55, n56, n57, n58, n59, n60, n61, n62, n63,
         n64, n65, n66, n67, n68, n69, n71, n74, n76, n77, n78, n79, n80, n81,
         n82, n83, n84, n86, n87, n88, n89, n90, n91, n92, n93, n94, n95, n96,
         n99, n100, n101, n102, n103, n105, n106, n107, n108, n109, n110, n111,
         n112, n113, n114, n115, n116, n117, n118, n119, n120, n122, n123,
         n124, n125, n126, n127, n128, n129, n130, n131, n132, n133, n134,
         n135, n136, n137, n139, n142, n144, n145, n146, n147, n148, n149,
         n150, n151, n152, n153, n154, n155, n156, n157, n158, n159, n160,
         n161, n162, n163, n164, n165, n166, n167, n169, n170, n171, n172,
         n173, n174, n176, n178, n179, n180, n181, n182, n187, n188, n189,
         n192, n194, n195, n196, n198, n200, n203, n205, n206, n207, n208,
         n209, n210, n211, n213, n215, n216, n217, n218, n219, n220, n222,
         n224, n225, n226, n228, n229, n230, n231, n233, n235, n236, n237,
         n240, n242, n243, n244, n245, n246, n248, n250, n252, n253, n254,
         n255, n256, n257, n258, n259, n260, n261, n262, n263, n264, n265,
         n266, n267, n268, n269, n270, n271, n272, n273, n275, n277, n278,
         n280, n282, n283, n284, n285, n286, n287, n288, n289, n290, n291,
         n292, n293, n294, n295, n297, n299, n300, n302, n304, n305, n306,
         n308, n310, n311, n312, n313, n314, n315, n316, n317, n318, n319,
         n320, n321, n322, n323, n324, n325, n326, n328, n330, n331, n332,
         n333, n334, n336, n338, n339, n340, n341, n343, n344, n346, n347,
         n348, n349, n350, n352, n354, n355, n356, n367, n369, n370, n373,
         n374, n378, n379, n380, n381, n383, n517, n518, n519, n520, n521,
         n522, n523, n524, n525, n526, n527, n528, n529, n530, n531, n532,
         n533, n534, n535, n536, n537, n538, n539, n540, n541, n542, n543,
         n544, n545, n546, n547, n548, n549, n550, n551;

  OAI21XL U433 ( .A0(n243), .A1(n237), .B0(n242), .Y(n236) );
  INVX3 U434 ( .A(n244), .Y(n243) );
  NOR2X2 U435 ( .A(B[7]), .B(A[7]), .Y(n312) );
  NAND2X1 U436 ( .A(B[36]), .B(A[39]), .Y(n79) );
  XOR2X1 U437 ( .A(n83), .B(n7), .Y(SUM[38]) );
  NAND2X2 U438 ( .A(B[32]), .B(A[32]), .Y(n136) );
  CLKBUFX3 U439 ( .A(n60), .Y(n517) );
  NOR2X2 U440 ( .A(n81), .B(n519), .Y(n76) );
  OR2X2 U441 ( .A(B[9]), .B(A[9]), .Y(n533) );
  NAND2X4 U442 ( .A(B[9]), .B(A[9]), .Y(n304) );
  NOR2X4 U443 ( .A(n149), .B(n146), .Y(n144) );
  OAI21X4 U444 ( .A0(n146), .A1(n150), .B0(n147), .Y(n145) );
  BUFX3 U445 ( .A(n158), .Y(n518) );
  NOR2X8 U446 ( .A(n110), .B(n117), .Y(n108) );
  NOR2X2 U447 ( .A(B[34]), .B(A[34]), .Y(n117) );
  BUFX4 U448 ( .A(n78), .Y(n519) );
  AOI21X1 U449 ( .A0(n527), .A1(n222), .B0(n213), .Y(n211) );
  INVX3 U450 ( .A(n224), .Y(n222) );
  AOI21XL U451 ( .A0(n145), .A1(n133), .B0(n134), .Y(n132) );
  AOI21X4 U452 ( .A0(n145), .A1(n126), .B0(n127), .Y(n125) );
  OAI21X1 U453 ( .A0(n107), .A1(n99), .B0(n100), .Y(n96) );
  OAI21X2 U454 ( .A0(n196), .A1(n173), .B0(n174), .Y(n172) );
  NAND2X2 U455 ( .A(n528), .B(n524), .Y(n173) );
  NAND2X2 U456 ( .A(B[33]), .B(A[33]), .Y(n129) );
  NOR2X2 U457 ( .A(n317), .B(n320), .Y(n315) );
  NOR2X4 U458 ( .A(B[5]), .B(A[5]), .Y(n320) );
  CLKINVX4 U459 ( .A(n124), .Y(n122) );
  NAND2X2 U460 ( .A(n144), .B(n126), .Y(n124) );
  NAND2XL U461 ( .A(n379), .B(n318), .Y(n39) );
  OAI21X2 U462 ( .A0(n317), .A1(n321), .B0(n318), .Y(n316) );
  NAND2X1 U463 ( .A(B[6]), .B(A[6]), .Y(n318) );
  NAND2X1 U464 ( .A(B[35]), .B(A[35]), .Y(n111) );
  BUFX3 U465 ( .A(n91), .Y(n520) );
  NOR2X4 U466 ( .A(B[33]), .B(A[33]), .Y(n128) );
  CLKINVX1 U467 ( .A(n77), .Y(n71) );
  AOI21X2 U468 ( .A0(n77), .A1(n58), .B0(n59), .Y(n57) );
  OAI21X2 U469 ( .A0(n519), .A1(n82), .B0(n79), .Y(n77) );
  BUFX4 U470 ( .A(n68), .Y(n521) );
  BUFX8 U471 ( .A(n90), .Y(n522) );
  INVX3 U472 ( .A(n200), .Y(n198) );
  NOR2X4 U473 ( .A(n128), .B(n135), .Y(n126) );
  AOI21X2 U474 ( .A0(n155), .A1(n542), .B0(n156), .Y(n154) );
  NOR2XL U475 ( .A(n169), .B(n162), .Y(n160) );
  NAND2X2 U476 ( .A(B[11]), .B(A[11]), .Y(n291) );
  XNOR2X2 U477 ( .A(n48), .B(n2), .Y(SUM[43]) );
  OAI21X2 U478 ( .A0(n110), .A1(n118), .B0(n111), .Y(n109) );
  NOR2X1 U479 ( .A(n99), .B(n522), .Y(n88) );
  CLKINVX1 U480 ( .A(n178), .Y(n176) );
  NAND2X1 U481 ( .A(n538), .B(n529), .Y(n230) );
  NAND2X1 U482 ( .A(n252), .B(n530), .Y(n245) );
  CLKINVX1 U483 ( .A(n250), .Y(n248) );
  AOI21X1 U484 ( .A0(n311), .A1(n535), .B0(n308), .Y(n306) );
  OAI21X1 U485 ( .A0(n326), .A1(n324), .B0(n325), .Y(n323) );
  NOR2X1 U486 ( .A(n106), .B(n99), .Y(n95) );
  NAND2X1 U487 ( .A(n76), .B(n58), .Y(n56) );
  NAND2X1 U488 ( .A(B[8]), .B(A[8]), .Y(n310) );
  OAI21X1 U489 ( .A0(n314), .A1(n312), .B0(n313), .Y(n311) );
  NAND2X1 U490 ( .A(B[13]), .B(A[13]), .Y(n282) );
  OR2X1 U491 ( .A(B[20]), .B(A[20]), .Y(n538) );
  NAND2X1 U492 ( .A(B[23]), .B(A[23]), .Y(n215) );
  NOR2X1 U493 ( .A(B[4]), .B(A[4]), .Y(n324) );
  NAND2X1 U494 ( .A(B[3]), .B(A[3]), .Y(n330) );
  AOI21X1 U495 ( .A0(n534), .A1(n339), .B0(n336), .Y(n334) );
  NOR2X1 U496 ( .A(B[2]), .B(A[2]), .Y(n332) );
  NAND2X1 U497 ( .A(B[1]), .B(A[1]), .Y(n338) );
  NAND2X1 U498 ( .A(B[0]), .B(A[0]), .Y(n341) );
  NOR2X2 U499 ( .A(B[30]), .B(A[30]), .Y(n149) );
  NOR2X1 U500 ( .A(B[36]), .B(A[37]), .Y(n90) );
  AOI21X1 U501 ( .A0(n206), .A1(n189), .B0(n194), .Y(n188) );
  XNOR2X1 U502 ( .A(n69), .B(n5), .Y(SUM[40]) );
  AOI21X1 U503 ( .A0(n206), .A1(n160), .B0(n161), .Y(n159) );
  XNOR2X1 U504 ( .A(n206), .B(n21), .Y(SUM[24]) );
  AOI21X1 U505 ( .A0(n206), .A1(n167), .B0(n542), .Y(n166) );
  AOI21X1 U506 ( .A0(n206), .A1(n180), .B0(n181), .Y(n179) );
  XNOR2X1 U507 ( .A(n112), .B(n10), .Y(SUM[35]) );
  OAI21X1 U508 ( .A0(n151), .A1(n113), .B0(n114), .Y(n112) );
  OAI21XL U509 ( .A0(n292), .A1(n290), .B0(n291), .Y(n289) );
  XNOR2X1 U510 ( .A(n101), .B(n9), .Y(SUM[36]) );
  OAI21X1 U511 ( .A0(n151), .A1(n142), .B0(n139), .Y(n137) );
  INVX4 U512 ( .A(n152), .Y(n151) );
  NOR2X2 U513 ( .A(B[32]), .B(A[32]), .Y(n135) );
  XNOR2X1 U514 ( .A(n130), .B(n12), .Y(SUM[33]) );
  OAI21X1 U515 ( .A0(n151), .A1(n131), .B0(n132), .Y(n130) );
  OAI21X1 U516 ( .A0(n83), .A1(n63), .B0(n64), .Y(n62) );
  INVX8 U517 ( .A(n545), .Y(n83) );
  OAI21X1 U518 ( .A0(n151), .A1(n149), .B0(n150), .Y(n148) );
  NOR2X2 U519 ( .A(B[36]), .B(A[36]), .Y(n99) );
  OR2X6 U520 ( .A(B[25]), .B(A[25]), .Y(n523) );
  OR2X4 U521 ( .A(B[27]), .B(A[27]), .Y(n524) );
  OR2X1 U522 ( .A(B[10]), .B(A[10]), .Y(n525) );
  OR2X1 U523 ( .A(B[14]), .B(A[14]), .Y(n526) );
  OR2X1 U524 ( .A(B[23]), .B(A[23]), .Y(n527) );
  OR2X2 U525 ( .A(B[26]), .B(A[26]), .Y(n528) );
  OR2X2 U526 ( .A(B[21]), .B(A[21]), .Y(n529) );
  OR2X1 U527 ( .A(B[19]), .B(A[19]), .Y(n530) );
  OR2X2 U528 ( .A(B[24]), .B(A[24]), .Y(n531) );
  OR2X1 U529 ( .A(B[13]), .B(A[13]), .Y(n532) );
  OR2X1 U530 ( .A(B[1]), .B(A[1]), .Y(n534) );
  OR2X1 U531 ( .A(B[8]), .B(A[8]), .Y(n535) );
  OR2X1 U532 ( .A(B[3]), .B(A[3]), .Y(n536) );
  OR2X1 U533 ( .A(B[22]), .B(A[22]), .Y(n537) );
  BUFX4 U534 ( .A(n172), .Y(n542) );
  NOR2X1 U535 ( .A(B[17]), .B(A[17]), .Y(n259) );
  INVX3 U536 ( .A(n242), .Y(n240) );
  OR2X1 U537 ( .A(n83), .B(n81), .Y(n541) );
  OR2X1 U538 ( .A(n151), .B(n102), .Y(n539) );
  NAND2X2 U539 ( .A(n539), .B(n103), .Y(n101) );
  OR2X1 U540 ( .A(n83), .B(n56), .Y(n540) );
  NAND2X2 U541 ( .A(n540), .B(n57), .Y(n55) );
  XNOR2X4 U542 ( .A(n55), .B(n3), .Y(SUM[42]) );
  NAND2X2 U543 ( .A(n541), .B(n82), .Y(n80) );
  XNOR2X4 U544 ( .A(n80), .B(n6), .Y(SUM[39]) );
  NAND2XL U545 ( .A(n122), .B(n115), .Y(n113) );
  OAI21X2 U546 ( .A0(n151), .A1(n120), .B0(n125), .Y(n119) );
  INVXL U547 ( .A(n122), .Y(n120) );
  NAND2XL U548 ( .A(n133), .B(n136), .Y(n13) );
  INVXL U549 ( .A(n136), .Y(n134) );
  OAI21X2 U550 ( .A0(n128), .A1(n136), .B0(n129), .Y(n127) );
  OAI21X1 U551 ( .A0(n157), .A1(n165), .B0(n518), .Y(n156) );
  AOI21X4 U552 ( .A0(n263), .A1(n271), .B0(n264), .Y(n262) );
  OAI21X1 U553 ( .A0(n265), .A1(n269), .B0(n266), .Y(n264) );
  NAND2XL U554 ( .A(n538), .B(n242), .Y(n25) );
  NAND2X2 U555 ( .A(B[20]), .B(A[20]), .Y(n242) );
  NOR2X2 U556 ( .A(n173), .B(n195), .Y(n171) );
  NAND2X1 U557 ( .A(B[27]), .B(A[27]), .Y(n178) );
  OAI21X2 U558 ( .A0(n151), .A1(n93), .B0(n94), .Y(n92) );
  NAND2X1 U559 ( .A(B[17]), .B(A[17]), .Y(n260) );
  NAND2XL U560 ( .A(n524), .B(n178), .Y(n18) );
  OAI21X1 U561 ( .A0(n83), .A1(n550), .B0(n549), .Y(n48) );
  XNOR2X2 U562 ( .A(n119), .B(n11), .Y(SUM[34]) );
  OAI21X1 U563 ( .A0(n83), .A1(n74), .B0(n71), .Y(n69) );
  NOR2X4 U564 ( .A(B[16]), .B(A[16]), .Y(n265) );
  NAND2X1 U565 ( .A(B[16]), .B(A[16]), .Y(n266) );
  CLKAND2X6 U566 ( .A(n285), .B(n293), .Y(n543) );
  NOR2X6 U567 ( .A(n543), .B(n286), .Y(n284) );
  OAI21X2 U568 ( .A0(n306), .A1(n294), .B0(n295), .Y(n293) );
  OAI21X4 U569 ( .A0(n287), .A1(n291), .B0(n288), .Y(n286) );
  INVXL U570 ( .A(n284), .Y(n283) );
  INVX8 U571 ( .A(n207), .Y(n206) );
  AND2XL U572 ( .A(B[26]), .B(A[26]), .Y(n544) );
  NAND2X2 U573 ( .A(B[22]), .B(A[22]), .Y(n224) );
  NOR2X6 U574 ( .A(B[35]), .B(A[35]), .Y(n110) );
  NOR2X6 U575 ( .A(B[6]), .B(A[6]), .Y(n317) );
  NOR2X6 U576 ( .A(B[12]), .B(A[12]), .Y(n287) );
  NAND2X6 U577 ( .A(B[30]), .B(A[30]), .Y(n150) );
  NOR2X4 U578 ( .A(B[29]), .B(A[29]), .Y(n157) );
  NAND2X4 U579 ( .A(B[28]), .B(A[28]), .Y(n165) );
  NOR2X1 U580 ( .A(B[11]), .B(A[11]), .Y(n290) );
  NAND2XL U581 ( .A(B[29]), .B(A[29]), .Y(n158) );
  NAND2XL U582 ( .A(B[12]), .B(A[12]), .Y(n288) );
  NOR2X1 U583 ( .A(B[28]), .B(A[28]), .Y(n164) );
  NOR2X1 U584 ( .A(n230), .B(n210), .Y(n208) );
  AOI21X4 U585 ( .A0(n244), .A1(n208), .B0(n209), .Y(n207) );
  OAI21X1 U586 ( .A0(n231), .A1(n210), .B0(n211), .Y(n209) );
  AOI21X2 U587 ( .A0(n529), .A1(n240), .B0(n233), .Y(n231) );
  NAND2X1 U588 ( .A(n526), .B(n532), .Y(n272) );
  NAND2XL U589 ( .A(n529), .B(n235), .Y(n24) );
  OA21X2 U590 ( .A0(n125), .A1(n86), .B0(n87), .Y(n546) );
  AOI21X1 U591 ( .A0(n524), .A1(n544), .B0(n176), .Y(n174) );
  CLKINVX3 U592 ( .A(n235), .Y(n233) );
  NAND2X1 U593 ( .A(B[36]), .B(A[38]), .Y(n82) );
  XOR2XL U594 ( .A(n151), .B(n15), .Y(SUM[30]) );
  NAND2X1 U595 ( .A(n525), .B(n533), .Y(n294) );
  INVXL U596 ( .A(n171), .Y(n169) );
  INVXL U597 ( .A(n542), .Y(n170) );
  INVXL U598 ( .A(n81), .Y(n347) );
  INVX3 U599 ( .A(n277), .Y(n275) );
  OAI21X1 U600 ( .A0(n170), .A1(n162), .B0(n165), .Y(n161) );
  INVX3 U601 ( .A(n299), .Y(n297) );
  OA21XL U602 ( .A0(n57), .A1(n53), .B0(n54), .Y(n549) );
  INVXL U603 ( .A(n254), .Y(n367) );
  OR2XL U604 ( .A(n56), .B(n53), .Y(n550) );
  OAI21XL U605 ( .A0(n270), .A1(n268), .B0(n269), .Y(n267) );
  OAI21XL U606 ( .A0(n322), .A1(n320), .B0(n321), .Y(n319) );
  INVX1 U607 ( .A(n195), .Y(n189) );
  INVX1 U608 ( .A(n228), .Y(n226) );
  INVXL U609 ( .A(n107), .Y(n105) );
  INVXL U610 ( .A(n145), .Y(n139) );
  NAND2X2 U611 ( .A(n531), .B(n523), .Y(n195) );
  OAI2BB1X4 U612 ( .A0N(n152), .A1N(n84), .B0(n546), .Y(n545) );
  OAI21X1 U613 ( .A0(n192), .A1(n182), .B0(n187), .Y(n181) );
  INVXL U614 ( .A(n528), .Y(n182) );
  INVXL U615 ( .A(n538), .Y(n237) );
  OAI21X4 U616 ( .A0(n153), .A1(n207), .B0(n154), .Y(n152) );
  NAND2X2 U617 ( .A(n155), .B(n171), .Y(n153) );
  OAI21X4 U618 ( .A0(n262), .A1(n245), .B0(n246), .Y(n244) );
  OAI21X4 U619 ( .A0(n284), .A1(n272), .B0(n273), .Y(n271) );
  AOI21X2 U620 ( .A0(n523), .A1(n203), .B0(n198), .Y(n196) );
  NAND2XL U621 ( .A(n349), .B(n100), .Y(n9) );
  INVXL U622 ( .A(n99), .Y(n349) );
  NAND2XL U623 ( .A(n354), .B(n147), .Y(n14) );
  OAI21X2 U624 ( .A0(n254), .A1(n260), .B0(n255), .Y(n253) );
  XNOR2X1 U625 ( .A(n547), .B(n20), .Y(SUM[25]) );
  AO21XL U626 ( .A0(n206), .A1(n531), .B0(n203), .Y(n547) );
  INVXL U627 ( .A(n522), .Y(n348) );
  INVXL U628 ( .A(n118), .Y(n116) );
  OAI21X2 U629 ( .A0(n334), .A1(n332), .B0(n333), .Y(n331) );
  XOR2XL U630 ( .A(n243), .B(n25), .Y(SUM[20]) );
  XNOR2X1 U631 ( .A(n548), .B(n26), .Y(SUM[19]) );
  AO21XL U632 ( .A0(n261), .A1(n252), .B0(n253), .Y(n548) );
  NAND2XL U633 ( .A(n367), .B(n255), .Y(n27) );
  INVXL U634 ( .A(n117), .Y(n115) );
  NAND2XL U635 ( .A(n526), .B(n277), .Y(n31) );
  AOI21XL U636 ( .A0(n283), .A1(n532), .B0(n280), .Y(n278) );
  XNOR2XL U637 ( .A(n261), .B(n28), .Y(SUM[17]) );
  XOR2XL U638 ( .A(n292), .B(n34), .Y(SUM[11]) );
  NAND2XL U639 ( .A(n525), .B(n299), .Y(n35) );
  AOI21XL U640 ( .A0(n305), .A1(n533), .B0(n302), .Y(n300) );
  XNOR2XL U641 ( .A(n283), .B(n32), .Y(SUM[13]) );
  XNOR2XL U642 ( .A(n305), .B(n36), .Y(SUM[9]) );
  XNOR2XL U643 ( .A(n311), .B(n37), .Y(SUM[8]) );
  XOR2XL U644 ( .A(n314), .B(n38), .Y(SUM[7]) );
  NAND2XL U645 ( .A(n378), .B(n313), .Y(n38) );
  INVXL U646 ( .A(n312), .Y(n378) );
  XOR2XL U647 ( .A(n41), .B(n326), .Y(SUM[4]) );
  NAND2XL U648 ( .A(n381), .B(n325), .Y(n41) );
  INVXL U649 ( .A(n324), .Y(n381) );
  XOR2XL U650 ( .A(n43), .B(n334), .Y(SUM[2]) );
  NAND2XL U651 ( .A(n383), .B(n333), .Y(n43) );
  INVXL U652 ( .A(n332), .Y(n383) );
  XNOR2XL U653 ( .A(n42), .B(n331), .Y(SUM[3]) );
  XNOR2XL U654 ( .A(n44), .B(n339), .Y(SUM[1]) );
  NOR2X4 U655 ( .A(B[31]), .B(A[31]), .Y(n146) );
  NAND2X2 U656 ( .A(B[24]), .B(A[24]), .Y(n205) );
  NAND2XL U657 ( .A(B[36]), .B(A[43]), .Y(n47) );
  NAND2XL U658 ( .A(B[36]), .B(A[40]), .Y(n68) );
  NAND2X4 U659 ( .A(B[15]), .B(A[15]), .Y(n269) );
  NAND2X4 U660 ( .A(B[5]), .B(A[5]), .Y(n321) );
  NOR2X4 U661 ( .A(B[18]), .B(A[18]), .Y(n254) );
  NAND2XL U662 ( .A(B[26]), .B(A[26]), .Y(n187) );
  NOR2X1 U663 ( .A(B[15]), .B(A[15]), .Y(n268) );
  NAND2XL U664 ( .A(B[36]), .B(A[37]), .Y(n91) );
  NOR2X1 U665 ( .A(B[36]), .B(A[39]), .Y(n78) );
  NOR2X1 U666 ( .A(B[36]), .B(A[40]), .Y(n67) );
  NOR2X1 U667 ( .A(B[36]), .B(A[38]), .Y(n81) );
  NOR2X1 U668 ( .A(B[36]), .B(A[41]), .Y(n60) );
  NOR2X1 U669 ( .A(B[36]), .B(A[42]), .Y(n53) );
  NAND2XL U670 ( .A(B[36]), .B(A[41]), .Y(n61) );
  NAND2XL U671 ( .A(B[36]), .B(A[42]), .Y(n54) );
  OR2XL U672 ( .A(B[36]), .B(A[43]), .Y(n551) );
  NAND2BXL U673 ( .AN(n340), .B(n341), .Y(n45) );
  NOR2XL U674 ( .A(B[0]), .B(A[0]), .Y(n340) );
  CLKINVX1 U675 ( .A(n169), .Y(n167) );
  NAND2X1 U676 ( .A(n122), .B(n108), .Y(n102) );
  AOI21X1 U677 ( .A0(n123), .A1(n108), .B0(n105), .Y(n103) );
  NAND2X1 U678 ( .A(n95), .B(n122), .Y(n93) );
  CLKINVX1 U679 ( .A(n230), .Y(n228) );
  NOR2X1 U680 ( .A(n195), .B(n182), .Y(n180) );
  NAND2X1 U681 ( .A(n228), .B(n219), .Y(n217) );
  NAND2X1 U682 ( .A(n537), .B(n527), .Y(n210) );
  CLKINVX1 U683 ( .A(n125), .Y(n123) );
  NAND2X1 U684 ( .A(n108), .B(n88), .Y(n86) );
  NOR2X1 U685 ( .A(n124), .B(n86), .Y(n84) );
  NAND2X1 U686 ( .A(n76), .B(n65), .Y(n63) );
  CLKINVX1 U687 ( .A(n76), .Y(n74) );
  AOI21X1 U688 ( .A0(n229), .A1(n219), .B0(n222), .Y(n218) );
  CLKINVX1 U689 ( .A(n262), .Y(n261) );
  CLKINVX1 U690 ( .A(n108), .Y(n106) );
  CLKINVX1 U691 ( .A(n144), .Y(n142) );
  CLKINVX1 U692 ( .A(n109), .Y(n107) );
  CLKINVX1 U693 ( .A(n231), .Y(n229) );
  CLKINVX1 U694 ( .A(n271), .Y(n270) );
  CLKINVX1 U695 ( .A(n220), .Y(n219) );
  CLKINVX1 U696 ( .A(n537), .Y(n220) );
  CLKINVX1 U697 ( .A(n194), .Y(n192) );
  CLKINVX1 U698 ( .A(n196), .Y(n194) );
  NAND2X1 U699 ( .A(n144), .B(n133), .Y(n131) );
  CLKINVX1 U700 ( .A(n293), .Y(n292) );
  CLKINVX1 U701 ( .A(n306), .Y(n305) );
  CLKINVX1 U702 ( .A(n323), .Y(n322) );
  CLKINVX1 U703 ( .A(n310), .Y(n308) );
  NOR2X1 U704 ( .A(n287), .B(n290), .Y(n285) );
  NOR2X1 U705 ( .A(n265), .B(n268), .Y(n263) );
  AOI21X1 U706 ( .A0(n253), .A1(n530), .B0(n248), .Y(n246) );
  NOR2X1 U707 ( .A(n157), .B(n164), .Y(n155) );
  AOI21X1 U708 ( .A0(n525), .A1(n302), .B0(n297), .Y(n295) );
  AOI21X1 U709 ( .A0(n526), .A1(n280), .B0(n275), .Y(n273) );
  AOI21X1 U710 ( .A0(n315), .A1(n323), .B0(n316), .Y(n314) );
  OAI21XL U711 ( .A0(n517), .A1(n521), .B0(n61), .Y(n59) );
  NAND2X1 U712 ( .A(n115), .B(n118), .Y(n11) );
  XNOR2X1 U713 ( .A(n137), .B(n13), .Y(SUM[32]) );
  XNOR2X1 U714 ( .A(n92), .B(n8), .Y(SUM[37]) );
  NAND2X1 U715 ( .A(n348), .B(n520), .Y(n8) );
  NAND2X1 U716 ( .A(n352), .B(n129), .Y(n12) );
  CLKINVX1 U717 ( .A(n128), .Y(n352) );
  XNOR2X1 U718 ( .A(n148), .B(n14), .Y(SUM[31]) );
  CLKINVX1 U719 ( .A(n146), .Y(n354) );
  NAND2X1 U720 ( .A(n350), .B(n111), .Y(n10) );
  CLKINVX1 U721 ( .A(n110), .Y(n350) );
  NAND2X1 U722 ( .A(n65), .B(n521), .Y(n5) );
  NAND2X1 U723 ( .A(n343), .B(n54), .Y(n3) );
  CLKINVX1 U724 ( .A(n53), .Y(n343) );
  XNOR2X1 U725 ( .A(n62), .B(n4), .Y(SUM[41]) );
  NAND2X1 U726 ( .A(n344), .B(n61), .Y(n4) );
  CLKINVX1 U727 ( .A(n517), .Y(n344) );
  NAND2X1 U728 ( .A(n346), .B(n79), .Y(n6) );
  CLKINVX1 U729 ( .A(n519), .Y(n346) );
  AOI21X1 U730 ( .A0(n109), .A1(n88), .B0(n89), .Y(n87) );
  OAI21XL U731 ( .A0(n522), .A1(n100), .B0(n520), .Y(n89) );
  AOI21X1 U732 ( .A0(n77), .A1(n65), .B0(n66), .Y(n64) );
  CLKINVX1 U733 ( .A(n521), .Y(n66) );
  AOI21X1 U734 ( .A0(n123), .A1(n115), .B0(n116), .Y(n114) );
  CLKINVX1 U735 ( .A(n215), .Y(n213) );
  AOI21X1 U736 ( .A0(n123), .A1(n95), .B0(n96), .Y(n94) );
  NOR2X1 U737 ( .A(n254), .B(n259), .Y(n252) );
  NOR2X1 U738 ( .A(n67), .B(n517), .Y(n58) );
  CLKINVX1 U739 ( .A(n67), .Y(n65) );
  CLKINVX1 U740 ( .A(n205), .Y(n203) );
  CLKINVX1 U741 ( .A(n282), .Y(n280) );
  CLKINVX1 U742 ( .A(n304), .Y(n302) );
  NAND2X1 U743 ( .A(n347), .B(n82), .Y(n7) );
  XOR2X1 U744 ( .A(n159), .B(n16), .Y(SUM[29]) );
  NAND2X1 U745 ( .A(n356), .B(n518), .Y(n16) );
  CLKINVX1 U746 ( .A(n157), .Y(n356) );
  XOR2X1 U747 ( .A(n166), .B(n17), .Y(SUM[28]) );
  NAND2X1 U748 ( .A(n163), .B(n165), .Y(n17) );
  XOR2X1 U749 ( .A(n179), .B(n18), .Y(SUM[27]) );
  XOR2X1 U750 ( .A(n188), .B(n19), .Y(SUM[26]) );
  NAND2X1 U751 ( .A(n528), .B(n187), .Y(n19) );
  NAND2X1 U752 ( .A(n523), .B(n200), .Y(n20) );
  NAND2X1 U753 ( .A(n355), .B(n150), .Y(n15) );
  CLKINVX1 U754 ( .A(n149), .Y(n355) );
  CLKINVX1 U755 ( .A(n338), .Y(n336) );
  AOI21X1 U756 ( .A0(n331), .A1(n536), .B0(n328), .Y(n326) );
  CLKINVX1 U757 ( .A(n330), .Y(n328) );
  NAND2X1 U758 ( .A(n531), .B(n205), .Y(n21) );
  XNOR2X1 U759 ( .A(n216), .B(n22), .Y(SUM[23]) );
  NAND2X1 U760 ( .A(n527), .B(n215), .Y(n22) );
  OAI21XL U761 ( .A0(n243), .A1(n217), .B0(n218), .Y(n216) );
  XNOR2X1 U762 ( .A(n225), .B(n23), .Y(SUM[22]) );
  NAND2X1 U763 ( .A(n219), .B(n224), .Y(n23) );
  OAI21XL U764 ( .A0(n243), .A1(n226), .B0(n231), .Y(n225) );
  XNOR2X1 U765 ( .A(n236), .B(n24), .Y(SUM[21]) );
  NAND2X1 U766 ( .A(n257), .B(n260), .Y(n28) );
  XNOR2X1 U767 ( .A(n267), .B(n29), .Y(SUM[16]) );
  NAND2X1 U768 ( .A(n369), .B(n266), .Y(n29) );
  CLKINVX1 U769 ( .A(n265), .Y(n369) );
  CLKINVX1 U770 ( .A(n135), .Y(n133) );
  CLKINVX1 U771 ( .A(n163), .Y(n162) );
  CLKINVX1 U772 ( .A(n164), .Y(n163) );
  CLKINVX1 U773 ( .A(n341), .Y(n339) );
  CLKINVX1 U774 ( .A(n259), .Y(n257) );
  XOR2X1 U775 ( .A(n270), .B(n30), .Y(SUM[15]) );
  NAND2X1 U776 ( .A(n370), .B(n269), .Y(n30) );
  CLKINVX1 U777 ( .A(n268), .Y(n370) );
  XOR2X1 U778 ( .A(n256), .B(n27), .Y(SUM[18]) );
  AOI21X1 U779 ( .A0(n261), .A1(n257), .B0(n258), .Y(n256) );
  XOR2X1 U780 ( .A(n278), .B(n31), .Y(SUM[14]) );
  NAND2X1 U781 ( .A(n530), .B(n250), .Y(n26) );
  CLKINVX1 U782 ( .A(n260), .Y(n258) );
  NAND2X1 U783 ( .A(n532), .B(n282), .Y(n32) );
  XNOR2X1 U784 ( .A(n289), .B(n33), .Y(SUM[12]) );
  NAND2X1 U785 ( .A(n373), .B(n288), .Y(n33) );
  CLKINVX1 U786 ( .A(n287), .Y(n373) );
  NAND2X1 U787 ( .A(n533), .B(n304), .Y(n36) );
  NAND2X1 U788 ( .A(n374), .B(n291), .Y(n34) );
  CLKINVX1 U789 ( .A(n290), .Y(n374) );
  XOR2X1 U790 ( .A(n300), .B(n35), .Y(SUM[10]) );
  XNOR2X1 U791 ( .A(n319), .B(n39), .Y(SUM[6]) );
  CLKINVX1 U792 ( .A(n317), .Y(n379) );
  NAND2X1 U793 ( .A(n535), .B(n310), .Y(n37) );
  XOR2X1 U794 ( .A(n40), .B(n322), .Y(SUM[5]) );
  NAND2X1 U795 ( .A(n380), .B(n321), .Y(n40) );
  CLKINVX1 U796 ( .A(n320), .Y(n380) );
  NAND2X1 U797 ( .A(n536), .B(n330), .Y(n42) );
  NAND2X1 U798 ( .A(n534), .B(n338), .Y(n44) );
  NAND2X1 U799 ( .A(n551), .B(n47), .Y(n2) );
  NAND2X1 U800 ( .A(B[34]), .B(A[34]), .Y(n118) );
  NAND2X1 U801 ( .A(B[36]), .B(A[36]), .Y(n100) );
  NAND2X1 U802 ( .A(B[25]), .B(A[25]), .Y(n200) );
  NAND2X1 U803 ( .A(B[21]), .B(A[21]), .Y(n235) );
  NAND2X1 U804 ( .A(B[14]), .B(A[14]), .Y(n277) );
  NAND2X1 U805 ( .A(B[10]), .B(A[10]), .Y(n299) );
  NAND2X1 U806 ( .A(B[19]), .B(A[19]), .Y(n250) );
  NAND2X1 U807 ( .A(B[31]), .B(A[31]), .Y(n147) );
  NAND2X1 U808 ( .A(B[18]), .B(A[18]), .Y(n255) );
  NAND2X1 U809 ( .A(B[4]), .B(A[4]), .Y(n325) );
  NAND2X1 U810 ( .A(B[7]), .B(A[7]), .Y(n313) );
  NAND2X1 U811 ( .A(B[2]), .B(A[2]), .Y(n333) );
  CLKINVX1 U812 ( .A(n45), .Y(SUM[0]) );
endmodule


module CONV ( clk, reset, busy, ready, iaddr, idata, cwr, caddr_wr, cdata_wr, 
        crd, caddr_rd, cdata_rd, csel );
  output [11:0] iaddr;
  input [19:0] idata;
  output [11:0] caddr_wr;
  output [19:0] cdata_wr;
  output [11:0] caddr_rd;
  input [19:0] cdata_rd;
  output [2:0] csel;
  input clk, reset, ready;
  output busy, cwr, crd;
  wire   n1132, n1133, n1134, n1135, n1136, n1137, n1138, n1139, n1140, n1141,
         n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, n1151,
         n1152, n1153, n1154, n1155, n1156, n1157, n1158, n1159, n1160,
         BiasTemp_7, N279, N281, N282, N283, N284, N314, N316, N317, N318,
         N319, N422, N430, N555, N556, N557, N558, N559, N560, N561, N562,
         N563, N564, N610, mulTemp_43, N703, N704, N705, N706, N707, N708,
         N709, N710, N711, N712, N713, N714, N715, N716, N717, N718, N719,
         N720, N721, N722, N723, N724, N725, N726, N727, N728, N729, N730,
         N731, N732, N733, N734, N735, N736, N737, N738, N739, N740, N741,
         N742, N743, N744, N745, N746, N1064, N1065, N1066, N1067, N1068,
         N1069, N1070, N1071, N1072, N1073, N1074, N1075, N1076, N1077, N1078,
         N1079, N1080, N1081, N1082, N1083, N1084, N1085, N1086, N1087, N1088,
         N1089, N1090, N1091, N1092, N1093, N1094, N1095, N1096, N1097, N1098,
         N1099, N1100, N1101, N1102, N1103, N1104, N1105, N1106, N1107, n28,
         n35, n36, n37, n38, n39, n40, n43, n44, n45, n46, n47, n78, n79, n80,
         n81, n92, n98, n99, n101, n117, n118, n120, n138, n142, n184, n185,
         n191, n192, n194, n198, n201, n202, n203, n204, n205, n206, n207,
         n209, n210, n211, n212, n213, n214, n235, n236, n262, n264, n265,
         n269, n277, n278, n279, n281, n282, n283, n284, n285, n286, n287,
         n289, n290, n291, n292, n293, n294, n296, n351, n359, n360, n367,
         n368, n369, n370, n371, n372, n373, n374, n375, n376, n377, n378,
         n379, n380, n381, n382, n383, n384, n385, n386, n387, n388, n389,
         n390, n391, n392, n393, n394, n395, n396, n397, n398, n399, n400,
         n401, n402, n403, n404, n405, n406, n407, n408, n409, n410, n411,
         n412, n413, n414, n415, n416, n417, n418, n419, n420, n421, n422,
         n423, n424, n425, n426, n427, n428, n429, n430, n431, n432, n433,
         n434, n435, n436, n437, n438, n439, n440, n441, n442, n443, n444,
         n445, n446, n447, n448, n449, n450, n451, n452, n453, n454, n455,
         n456, n457, n458, n459, n460, n461, n462, n463, n464, n465, n466,
         n467, n468, \add_153_S2/carry[5] , \add_153_S2/carry[4] ,
         \add_153_S2/carry[3] , \add_140/carry[5] , \add_140/carry[4] ,
         \add_140/carry[3] , \r363/carry[5] , \r363/carry[4] , \r363/carry[3] ,
         \r363/carry[2] , \r361/carry[5] , \r361/carry[4] , \r361/carry[3] ,
         \r361/carry[2] , n469, n470, n471, n472, n473, n474, n475, n476, n477,
         n478, n479, n480, n481, n482, n483, n484, n485, n486, n487, n488,
         n489, n490, n491, n492, n493, n494, n495, n496, n497, n498, n500,
         n502, n503, n504, n505, n506, n507, n508, n509, n510, n511, n512,
         n513, n514, n515, n516, n517, n518, n519, n520, n521, n522, n523,
         n524, n525, n526, n527, n528, n529, n530, n531, n532, n533, n534,
         n535, n536, n537, n538, n539, n540, n541, n542, n543, n544, n545,
         n546, n547, n548, n549, n550, n551, n552, n553, n554, n555, n556,
         n557, n558, n559, n560, n561, n562, n564, n566, n568, n570, n572,
         n574, n578, n580, n582, n584, n1163, n586, n588, n590, n592, n594,
         n596, n598, n600, n602, n604, n606, n608, n610, n612, n614, n616,
         n618, n620, n622, n624, n626, n628, n630, n632, n634, n636, n638,
         n640, n642, n644, n646, n648, n650, n652, n654, n656, n658, n660,
         n662, n664, n666, n668, n670, n672, n674, n676, n678, n680, n682,
         n683, n684, n685, n686, n687, n688, n689, n690, n691, n692, n693,
         n694, n695, n696, n697, n698, n699, n700, n701, n702, n703, n704,
         n705, n706, n707, n708, n709, n710, n711, n712, n713, n714, n715,
         n716, n717, n718, n719, n720, n721, n722, n723, n724, n725, n726,
         n727, n728, n729, n730, n731, n732, n733, n734, n735, n736, n737,
         n738, n739, n740, n741, n742, n743, n744, n745, n746, n747, n748,
         n749, n750, n751, n752, n753, n754, n755, n756, n757, n758, n759,
         n760, n761, n762, n763, n764, n765, n766, n767, n768, n769, n770,
         n771, n772, n773, n774, n775, n776, n777, n778, n779, n780, n781,
         n782, n783, n784, n785, n786, n787, n788, n789, n790, n791, n792,
         n793, n794, n795, n796, n797, n798, n799, n800, n801, n802, n803,
         n804, n805, n806, n807, n808, n809, n810, n811, n812, n813, n814,
         n815, n816, n817, n818, n819, n820, n821, n822, n823, n824, n825,
         n826, n827, n828, n829, n830, n831, n832, n833, n834, n835, n836,
         n837, n838, n839, n840, n841, n842, n843, n844, n845, n846, n847,
         n848, n849, n850, n851, n852, n853, n854, n855, n856, n857, n858,
         n859, n860, n861, n862, n863, n864, n865, n866, n867, n868, n869,
         n870, n871, n872, n873, n874, n875, n876, n877, n878, n879, n880,
         n881, n882, n883, n884, n885, n886, n887, n888, n889, n890, n891,
         n892, n893, n894, n895, n896, n897, n898, n899, n900, n901, n902,
         n903, n904, n905, n906, n907, n908, n909, n910, n911, n912, n913,
         n914, n915, n916, n917, n918, n919, n920, n921, n922, n923, n924,
         n925, n926, n927, n928, n929, n930, n931, n932, n933, n934, n935,
         n936, n937, n938, n939, n940, n941, n942, n943, n944, n945, n946,
         n947, n948, n949, n950, n951, n952, n953, n954, n955, n956, n957,
         n958, n959, n960, n961, n962, n963, n964, n965, n966, n967, n968,
         n969, n970, n971, n972, n973, n974, n975, n976, n977, n978, n979,
         n980, n981, n982, n983, n984, n985, n986, n987, n988, n989, n990,
         n991, n992, n993, n994, n995, n996, n997, n998, n999, n1000, n1001,
         n1002, n1003, n1004, n1005, n1006, n1007, n1008, n1009, n1010, n1011,
         n1012, n1013, n1014, n1015, n1016, n1017, n1018, n1019, n1020, n1021,
         n1022, n1023, n1024, n1025, n1026, n1027, n1028, n1029, n1030, n1031,
         n1032, n1033, n1034, n1035, n1036, n1037, n1038, n1039, n1040, n1041,
         n1042, n1043, n1044, n1045, n1046, n1047, n1048, n1049, n1050, n1051,
         n1052, n1053, n1054, n1055, n1056, n1057, n1058, n1059, n1060, n1061,
         n1062, n1063, n1064, n1065, n1066, n1067, n1068, n1069, n1070, n1071,
         n1072, n1073, n1074, n1075, n1076, n1077, n1078, n1079, n1080, n1081,
         n1082, n1083, n1084, n1085, n1086, n1087, n1088, n1089, n1090, n1091,
         n1092, n1093, n1094, n1095, n1096, n1097, n1098, n1099, n1100, n1101,
         n1102, n1103, n1104, n1105, n1106, n1107, n1108, n1109, n1110, n1111,
         n1112, n1113, n1114, n1115, n1116, n1117, n1118, n1119, n1120, n1121,
         n1122, n1123, n1124, n1125, n1126, n1127, n1128, n1129, n1130, n1131,
         n1161;
  wire   [43:0] convTemp;
  wire   [20:1] roundTemp;
  wire   [3:0] counterRead;
  wire   [3:0] current_State;
  wire   [19:0] kernelTemp;
  wire   [5:0] index_X_Before;
  wire   [5:0] index_X_After;
  wire   [5:0] index_Y_Before;
  wire   [5:0] index_Y_After;
  wire   [3:0] next_State;
  wire   [19:0] idataTemp;
  wire   [38:0] mulTemp;
  wire   SYNOPSYS_UNCONNECTED__0;

  DFFRX1 \index_Y_reg[5]  ( .D(n464), .CK(clk), .RN(n740), .Q(N564), .QN(n40)
         );
  DFFRX1 \index_Y_reg[4]  ( .D(n458), .CK(clk), .RN(n740), .Q(N563), .QN(n43)
         );
  DFFRX1 \index_Y_reg[3]  ( .D(n459), .CK(clk), .RN(n739), .Q(N562), .QN(n44)
         );
  DFFRX2 \index_X_reg[1]  ( .D(n456), .CK(clk), .RN(n740), .Q(N555), .QN(n38)
         );
  DFFRX2 \index_X_reg[2]  ( .D(n455), .CK(clk), .RN(n740), .Q(N556), .QN(n37)
         );
  DFFRX2 \index_Y_reg[0]  ( .D(n462), .CK(clk), .RN(n740), .Q(N314), .QN(n47)
         );
  DFFRX2 \index_X_reg[0]  ( .D(n457), .CK(clk), .RN(n740), .Q(N279), .QN(n39)
         );
  EDFFX1 \idataTemp_reg[18]  ( .D(idata[18]), .E(n495), .CK(clk), .Q(
        idataTemp[18]) );
  EDFFX1 \idataTemp_reg[14]  ( .D(idata[14]), .E(n495), .CK(clk), .Q(
        idataTemp[14]) );
  EDFFX1 \idataTemp_reg[10]  ( .D(idata[10]), .E(n495), .CK(clk), .Q(
        idataTemp[10]) );
  EDFFX1 \idataTemp_reg[8]  ( .D(idata[8]), .E(n495), .CK(clk), .Q(
        idataTemp[8]) );
  EDFFX1 \idataTemp_reg[4]  ( .D(idata[4]), .E(n495), .CK(clk), .Q(
        idataTemp[4]) );
  EDFFX1 \idataTemp_reg[2]  ( .D(idata[2]), .E(n495), .CK(clk), .Q(
        idataTemp[2]) );
  EDFFX1 \idataTemp_reg[17]  ( .D(idata[17]), .E(n495), .CK(clk), .Q(
        idataTemp[17]) );
  EDFFX1 \idataTemp_reg[15]  ( .D(idata[15]), .E(n495), .CK(clk), .Q(
        idataTemp[15]) );
  EDFFX1 \idataTemp_reg[13]  ( .D(idata[13]), .E(n495), .CK(clk), .Q(
        idataTemp[13]) );
  EDFFX1 \idataTemp_reg[11]  ( .D(idata[11]), .E(n495), .CK(clk), .Q(
        idataTemp[11]) );
  EDFFX1 \idataTemp_reg[9]  ( .D(idata[9]), .E(n495), .CK(clk), .Q(
        idataTemp[9]) );
  EDFFX1 \idataTemp_reg[7]  ( .D(idata[7]), .E(n495), .CK(clk), .Q(
        idataTemp[7]) );
  EDFFX1 \idataTemp_reg[5]  ( .D(idata[5]), .E(n495), .CK(clk), .Q(
        idataTemp[5]) );
  EDFFX1 \idataTemp_reg[3]  ( .D(idata[3]), .E(n495), .CK(clk), .Q(
        idataTemp[3]) );
  EDFFX1 \idataTemp_reg[1]  ( .D(idata[1]), .E(n495), .CK(clk), .Q(
        idataTemp[1]) );
  EDFFX1 \idataTemp_reg[0]  ( .D(idata[0]), .E(n495), .CK(clk), .Q(
        idataTemp[0]) );
  DFFRX1 \convTemp_reg[43]  ( .D(n369), .CK(clk), .RN(n737), .Q(convTemp[43])
         );
  DFFRX1 \convTemp_reg[36]  ( .D(n376), .CK(clk), .RN(n736), .Q(convTemp[36]), 
        .QN(n1032) );
  DFFRX1 \convTemp_reg[37]  ( .D(n375), .CK(clk), .RN(n736), .Q(convTemp[37]), 
        .QN(n1028) );
  DFFRX1 \index_X_reg[4]  ( .D(n453), .CK(clk), .RN(n740), .Q(N558), .QN(n35)
         );
  DFFRX1 \index_X_reg[3]  ( .D(n454), .CK(clk), .RN(n740), .Q(N557), .QN(n36)
         );
  DFFRX1 \convTemp_reg[7]  ( .D(n406), .CK(clk), .RN(n734), .Q(convTemp[7]), 
        .QN(n967) );
  DFFRX1 \convTemp_reg[10]  ( .D(n403), .CK(clk), .RN(n734), .Q(convTemp[10]), 
        .QN(n955) );
  DFFRX1 \convTemp_reg[12]  ( .D(n401), .CK(clk), .RN(n734), .Q(convTemp[12]), 
        .QN(n947) );
  DFFRX1 \convTemp_reg[14]  ( .D(n399), .CK(clk), .RN(n734), .Q(convTemp[14]), 
        .QN(n939) );
  DFFRX1 \index_Y_reg[2]  ( .D(n460), .CK(clk), .RN(n740), .Q(N561), .QN(n45)
         );
  DFFRX1 \convTemp_reg[35]  ( .D(n378), .CK(clk), .RN(n735), .Q(convTemp[35]), 
        .QN(n1003) );
  DFFRX1 \index_Y_reg[1]  ( .D(n461), .CK(clk), .RN(n740), .Q(N560), .QN(n46)
         );
  DFFRX1 \convTemp_reg[33]  ( .D(n380), .CK(clk), .RN(n732), .Q(convTemp[33]), 
        .QN(n863) );
  DFFRX1 \convTemp_reg[34]  ( .D(n379), .CK(clk), .RN(n735), .Q(convTemp[34]), 
        .QN(n999) );
  DFFRX1 \convTemp_reg[31]  ( .D(n382), .CK(clk), .RN(n732), .Q(convTemp[31]), 
        .QN(n871) );
  DFFRX1 \convTemp_reg[0]  ( .D(n413), .CK(clk), .RN(n735), .Q(convTemp[0]), 
        .QN(n995) );
  DFFRX1 \convTemp_reg[1]  ( .D(n412), .CK(clk), .RN(n735), .Q(convTemp[1]), 
        .QN(n991) );
  DFFRX1 \convTemp_reg[2]  ( .D(n411), .CK(clk), .RN(n735), .Q(convTemp[2]), 
        .QN(n987) );
  DFFRX1 \convTemp_reg[3]  ( .D(n410), .CK(clk), .RN(n735), .Q(convTemp[3]), 
        .QN(n983) );
  DFFRX1 \convTemp_reg[4]  ( .D(n409), .CK(clk), .RN(n735), .Q(convTemp[4]), 
        .QN(n979) );
  DFFRX1 \convTemp_reg[5]  ( .D(n408), .CK(clk), .RN(n735), .Q(convTemp[5]), 
        .QN(n975) );
  DFFRX1 \convTemp_reg[6]  ( .D(n407), .CK(clk), .RN(n734), .Q(convTemp[6]), 
        .QN(n971) );
  DFFRX1 \convTemp_reg[27]  ( .D(n386), .CK(clk), .RN(n733), .Q(convTemp[27]), 
        .QN(n887) );
  DFFRX1 \convTemp_reg[25]  ( .D(n388), .CK(clk), .RN(n733), .Q(convTemp[25]), 
        .QN(n895) );
  DFFRX1 \convTemp_reg[23]  ( .D(n390), .CK(clk), .RN(n733), .Q(convTemp[23]), 
        .QN(n903) );
  DFFRX1 \convTemp_reg[21]  ( .D(n392), .CK(clk), .RN(n733), .Q(convTemp[21]), 
        .QN(n911) );
  DFFRX1 \convTemp_reg[22]  ( .D(n391), .CK(clk), .RN(n733), .Q(convTemp[22]), 
        .QN(n907) );
  DFFRX4 \counterRead_reg[3]  ( .D(n467), .CK(clk), .RN(n732), .Q(
        counterRead[3]), .QN(n92) );
  DFFRX4 \counterRead_reg[2]  ( .D(n465), .CK(clk), .RN(n732), .Q(
        counterRead[2]), .QN(n98) );
  DFFRX1 \convTemp_reg[20]  ( .D(n393), .CK(clk), .RN(n733), .Q(convTemp[20]), 
        .QN(n915) );
  DFFRX1 \convTemp_reg[19]  ( .D(n394), .CK(clk), .RN(n733), .Q(convTemp[19]), 
        .QN(n919) );
  DFFRX1 \convTemp_reg[13]  ( .D(n400), .CK(clk), .RN(n734), .Q(convTemp[13]), 
        .QN(n943) );
  DFFRX1 \convTemp_reg[8]  ( .D(n405), .CK(clk), .RN(n734), .Q(convTemp[8]), 
        .QN(n963) );
  DFFRX1 \convTemp_reg[9]  ( .D(n404), .CK(clk), .RN(n734), .Q(convTemp[9]), 
        .QN(n959) );
  DFFRX1 \convTemp_reg[11]  ( .D(n402), .CK(clk), .RN(n734), .Q(convTemp[11]), 
        .QN(n951) );
  DFFRX1 \convTemp_reg[32]  ( .D(n381), .CK(clk), .RN(n732), .Q(convTemp[32]), 
        .QN(n867) );
  DFFRX1 \convTemp_reg[30]  ( .D(n383), .CK(clk), .RN(n732), .Q(convTemp[30]), 
        .QN(n875) );
  DFFRX1 \convTemp_reg[24]  ( .D(n389), .CK(clk), .RN(n733), .Q(convTemp[24]), 
        .QN(n899) );
  DFFRX4 \counterRead_reg[0]  ( .D(n468), .CK(clk), .RN(n732), .Q(
        counterRead[0]), .QN(n101) );
  DFFRX1 \convTemp_reg[29]  ( .D(n384), .CK(clk), .RN(n733), .Q(convTemp[29]), 
        .QN(n879) );
  DFFRX4 \counterRead_reg[1]  ( .D(n466), .CK(clk), .RN(n732), .Q(
        counterRead[1]), .QN(n99) );
  DFFRX1 \convTemp_reg[42]  ( .D(n370), .CK(clk), .RN(n735), .Q(convTemp[42]), 
        .QN(n1011) );
  DFFRX1 \convTemp_reg[40]  ( .D(n372), .CK(clk), .RN(n735), .Q(convTemp[40]), 
        .QN(n1017) );
  DFFRX1 \convTemp_reg[38]  ( .D(n374), .CK(clk), .RN(n736), .Q(convTemp[38]), 
        .QN(n1024) );
  DFFRX1 \convTemp_reg[39]  ( .D(n373), .CK(clk), .RN(n735), .Q(convTemp[39]), 
        .QN(n1020) );
  DFFRX1 \convTemp_reg[15]  ( .D(n398), .CK(clk), .RN(n734), .Q(convTemp[15]), 
        .QN(n935) );
  DFFRX1 \convTemp_reg[17]  ( .D(n396), .CK(clk), .RN(n734), .Q(convTemp[17]), 
        .QN(n927) );
  DFFRX4 \current_State_reg[2]  ( .D(next_State[2]), .CK(clk), .RN(n732), .Q(
        current_State[2]), .QN(n79) );
  DFFRX1 \caddr_wr_reg[11]  ( .D(n474), .CK(clk), .RN(n738), .Q(n1135), .QN(
        n654) );
  DFFRX1 \csel_reg[0]  ( .D(n449), .CK(clk), .RN(n739), .Q(n1160), .QN(n652)
         );
  DFFRX1 \csel_reg[2]  ( .D(n451), .CK(clk), .RN(n739), .Q(n1158), .QN(n650)
         );
  DFFRX1 \csel_reg[1]  ( .D(n450), .CK(clk), .RN(n739), .Q(n1159), .QN(n648)
         );
  DFFRX1 \caddr_rd_reg[10]  ( .D(n435), .CK(clk), .RN(n739), .Q(n1157), .QN(
        n646) );
  DFFRX1 \caddr_rd_reg[11]  ( .D(n436), .CK(clk), .RN(n739), .Q(n1156), .QN(
        n644) );
  DFFRX1 \caddr_wr_reg[0]  ( .D(n414), .CK(clk), .RN(n738), .QN(n642) );
  DFFRX1 \iaddr_reg[4]  ( .D(n441), .CK(clk), .RN(n741), .QN(n640) );
  DFFRX1 \iaddr_reg[5]  ( .D(n442), .CK(clk), .RN(n741), .QN(n638) );
  DFFRX1 \iaddr_reg[10]  ( .D(n447), .CK(clk), .RN(n742), .QN(n636) );
  DFFRX1 \iaddr_reg[11]  ( .D(n448), .CK(clk), .RN(n742), .QN(n634) );
  DFFRX1 \caddr_wr_reg[6]  ( .D(n420), .CK(clk), .RN(n738), .QN(n632) );
  DFFRX1 \caddr_wr_reg[7]  ( .D(n421), .CK(clk), .RN(n738), .QN(n630) );
  DFFRX1 \caddr_wr_reg[8]  ( .D(n422), .CK(clk), .RN(n738), .QN(n628) );
  DFFRX1 \caddr_wr_reg[9]  ( .D(n423), .CK(clk), .RN(n738), .QN(n626) );
  DFFRX1 \iaddr_reg[3]  ( .D(n440), .CK(clk), .RN(n741), .QN(n624) );
  DFFRX1 \iaddr_reg[9]  ( .D(n446), .CK(clk), .RN(n742), .QN(n622) );
  DFFRX1 \caddr_wr_reg[1]  ( .D(n415), .CK(clk), .RN(n738), .QN(n620) );
  DFFRX1 \caddr_wr_reg[2]  ( .D(n416), .CK(clk), .RN(n738), .QN(n618) );
  DFFRX1 \caddr_wr_reg[3]  ( .D(n417), .CK(clk), .RN(n738), .QN(n616) );
  DFFRX1 \caddr_wr_reg[4]  ( .D(n418), .CK(clk), .RN(n738), .QN(n614) );
  DFFRX1 \caddr_wr_reg[5]  ( .D(n419), .CK(clk), .RN(n738), .QN(n612) );
  DFFRX1 \caddr_wr_reg[10]  ( .D(n424), .CK(clk), .RN(n741), .QN(n610) );
  DFFRX1 \caddr_rd_reg[0]  ( .D(n425), .CK(clk), .RN(n738), .QN(n608) );
  DFFRX1 \caddr_rd_reg[1]  ( .D(n426), .CK(clk), .RN(n739), .QN(n606) );
  DFFRX1 \caddr_rd_reg[2]  ( .D(n427), .CK(clk), .RN(n739), .QN(n604) );
  DFFRX1 \caddr_rd_reg[3]  ( .D(n428), .CK(clk), .RN(n739), .QN(n602) );
  DFFRX1 \caddr_rd_reg[4]  ( .D(n429), .CK(clk), .RN(n739), .QN(n600) );
  DFFRX1 \caddr_rd_reg[5]  ( .D(n430), .CK(clk), .RN(n739), .QN(n598) );
  DFFRX1 \caddr_rd_reg[6]  ( .D(n431), .CK(clk), .RN(n740), .QN(n596) );
  DFFRX1 \caddr_rd_reg[7]  ( .D(n432), .CK(clk), .RN(n741), .QN(n594) );
  DFFRX1 \caddr_rd_reg[8]  ( .D(n433), .CK(clk), .RN(n741), .QN(n592) );
  DFFRX1 \caddr_rd_reg[9]  ( .D(n434), .CK(clk), .RN(n741), .QN(n590) );
  DFFRX1 \iaddr_reg[1]  ( .D(n438), .CK(clk), .RN(n741), .QN(n588) );
  DFFRX1 \iaddr_reg[2]  ( .D(n439), .CK(clk), .RN(n741), .QN(n586) );
  DFFRX1 \iaddr_reg[8]  ( .D(n445), .CK(clk), .RN(n742), .QN(n582) );
  DFFRX1 busy_reg ( .D(n452), .CK(clk), .RN(n742), .Q(n1132), .QN(n580) );
  DFFRX1 \iaddr_reg[0]  ( .D(n437), .CK(clk), .RN(n741), .Q(n1134), .QN(n578)
         );
  DFFRX1 \iaddr_reg[6]  ( .D(n443), .CK(clk), .RN(n741), .Q(n1133), .QN(n702)
         );
  DFFRX1 cwr_reg ( .D(N422), .CK(clk), .RN(n739), .QN(n498) );
  DFFRX2 \current_State_reg[1]  ( .D(next_State[1]), .CK(clk), .RN(n732), .Q(
        current_State[1]), .QN(n80) );
  EDFFXL \idataTemp_reg[19]  ( .D(idata[19]), .E(n495), .CK(clk), .Q(
        idataTemp[19]) );
  EDFFXL \idataTemp_reg[16]  ( .D(idata[16]), .E(n495), .CK(clk), .Q(
        idataTemp[16]) );
  EDFFXL \idataTemp_reg[12]  ( .D(idata[12]), .E(n495), .CK(clk), .Q(
        idataTemp[12]) );
  EDFFXL \idataTemp_reg[6]  ( .D(idata[6]), .E(n495), .CK(clk), .Q(
        idataTemp[6]) );
  DFFRX4 \current_State_reg[3]  ( .D(next_State[3]), .CK(clk), .RN(n1112), .Q(
        current_State[3]), .QN(n78) );
  DFFRX1 \index_X_reg[5]  ( .D(n463), .CK(clk), .RN(n740), .Q(N559), .QN(n28)
         );
  DFFRX1 \cdata_wr_reg[0]  ( .D(n1122), .CK(clk), .RN(n737), .Q(n1155), .QN(
        n668) );
  DFFRX1 \convTemp_reg[28]  ( .D(n385), .CK(clk), .RN(n733), .Q(convTemp[28]), 
        .QN(n883) );
  DFFRX1 \convTemp_reg[26]  ( .D(n387), .CK(clk), .RN(n733), .Q(convTemp[26]), 
        .QN(n891) );
  DFFRX1 \convTemp_reg[41]  ( .D(n371), .CK(clk), .RN(n735), .Q(convTemp[41]), 
        .QN(n1014) );
  DFFRX1 \convTemp_reg[18]  ( .D(n395), .CK(clk), .RN(n733), .Q(convTemp[18]), 
        .QN(n923) );
  DFFRX1 \cdata_wr_reg[19]  ( .D(n377), .CK(clk), .RN(n737), .Q(n1136), .QN(
        n678) );
  DFFRX2 \current_State_reg[0]  ( .D(next_State[0]), .CK(clk), .RN(n732), .Q(
        current_State[0]), .QN(n81) );
  DFFRX1 \convTemp_reg[16]  ( .D(n397), .CK(clk), .RN(n734), .Q(convTemp[16]), 
        .QN(n931) );
  DFFRX1 \cdata_wr_reg[1]  ( .D(n492), .CK(clk), .RN(n736), .Q(n1154), .QN(
        n566) );
  DFFRX1 \cdata_wr_reg[2]  ( .D(n491), .CK(clk), .RN(n736), .Q(n1153), .QN(
        n568) );
  DFFRX1 \cdata_wr_reg[3]  ( .D(n490), .CK(clk), .RN(n736), .Q(n1152), .QN(
        n672) );
  DFFRX1 \cdata_wr_reg[4]  ( .D(n489), .CK(clk), .RN(n736), .Q(n1151), .QN(
        n664) );
  DFFRX1 \cdata_wr_reg[5]  ( .D(n488), .CK(clk), .RN(n736), .Q(n1150), .QN(
        n676) );
  DFFRX1 \cdata_wr_reg[6]  ( .D(n487), .CK(clk), .RN(n736), .Q(n1149), .QN(
        n658) );
  DFFRX1 \cdata_wr_reg[7]  ( .D(n486), .CK(clk), .RN(n736), .Q(n1148), .QN(
        n564) );
  DFFRX1 \cdata_wr_reg[8]  ( .D(n485), .CK(clk), .RN(n736), .Q(n1147), .QN(
        n674) );
  DFFRX1 \cdata_wr_reg[9]  ( .D(n484), .CK(clk), .RN(n736), .Q(n1146), .QN(
        n666) );
  DFFRX1 \cdata_wr_reg[10]  ( .D(n483), .CK(clk), .RN(n737), .Q(n1145), .QN(
        n570) );
  DFFRX1 \cdata_wr_reg[11]  ( .D(n482), .CK(clk), .RN(n737), .Q(n1144), .QN(
        n662) );
  DFFRX1 \cdata_wr_reg[12]  ( .D(n481), .CK(clk), .RN(n737), .Q(n1143), .QN(
        n680) );
  DFFRX1 \cdata_wr_reg[13]  ( .D(n480), .CK(clk), .RN(n737), .Q(n1142), .QN(
        n660) );
  DFFRX1 \cdata_wr_reg[14]  ( .D(n479), .CK(clk), .RN(n737), .Q(n1141), .QN(
        n572) );
  DFFRX1 \cdata_wr_reg[15]  ( .D(n478), .CK(clk), .RN(n737), .Q(n1140), .QN(
        n656) );
  DFFRX1 \cdata_wr_reg[16]  ( .D(n477), .CK(clk), .RN(n737), .Q(n1139), .QN(
        n562) );
  DFFRX1 \cdata_wr_reg[17]  ( .D(n476), .CK(clk), .RN(n737), .Q(n1138), .QN(
        n574) );
  DFFRX1 \cdata_wr_reg[18]  ( .D(n475), .CK(clk), .RN(n737), .Q(n1137), .QN(
        n670) );
  NAND3BX1 U460 ( .AN(n1023), .B(n1019), .C(n1018), .Y(n372) );
  AO21XL U461 ( .A0(n764), .A1(n776), .B0(current_State[3]), .Y(next_State[3])
         );
  OAI211XL U462 ( .A0(current_State[3]), .A1(n744), .B0(n1065), .C0(n853), .Y(
        n745) );
  NAND2XL U463 ( .A(n694), .B(current_State[3]), .Y(n782) );
  CLKINVX8 U464 ( .A(current_State[2]), .Y(n469) );
  INVX8 U465 ( .A(n469), .Y(n470) );
  INVX1 U466 ( .A(n469), .Y(n471) );
  NAND2X2 U467 ( .A(n1035), .B(n1034), .Y(n376) );
  AOI2BB2X2 U468 ( .B0(N739), .B1(n724), .A0N(n720), .A1N(n1027), .Y(n1035) );
  NOR3X8 U469 ( .A(n81), .B(n470), .C(current_State[3]), .Y(n685) );
  AND2X1 U470 ( .A(n471), .B(n78), .Y(n693) );
  NAND3BXL U471 ( .AN(n471), .B(n78), .C(n694), .Y(n788) );
  NOR2XL U472 ( .A(current_State[1]), .B(n471), .Y(n704) );
  NAND3BX2 U473 ( .AN(n1023), .B(n1022), .C(n1021), .Y(n373) );
  NAND2X2 U474 ( .A(N742), .B(n724), .Y(n1022) );
  AND2X6 U475 ( .A(n823), .B(n830), .Y(n687) );
  INVXL U476 ( .A(mulTemp[33]), .Y(n861) );
  AOI222X1 U477 ( .A0(n1155), .A1(n709), .B0(cdata_rd[0]), .B1(n710), .C0(
        roundTemp[1]), .C1(n711), .Y(n138) );
  BUFX12 U478 ( .A(n118), .Y(n710) );
  CLKBUFX8 U479 ( .A(n117), .Y(n709) );
  NAND3BX2 U480 ( .AN(n1023), .B(n1013), .C(n1012), .Y(n370) );
  AOI2BB2X2 U481 ( .B0(N1106), .B1(n686), .A0N(n722), .A1N(n1011), .Y(n1012)
         );
  AOI2BB2X4 U482 ( .B0(N1105), .B1(n727), .A0N(n722), .A1N(n1014), .Y(n1015)
         );
  NAND2X6 U483 ( .A(n101), .B(n1050), .Y(n1074) );
  NAND2X1 U484 ( .A(n806), .B(n805), .Y(n820) );
  NAND2X2 U485 ( .A(n692), .B(n843), .Y(n799) );
  NAND2X1 U486 ( .A(n813), .B(n1123), .Y(n814) );
  AO21X1 U487 ( .A0(n1050), .A1(n707), .B0(n700), .Y(n817) );
  NAND2X2 U488 ( .A(n1093), .B(n820), .Y(n815) );
  NAND2X1 U489 ( .A(n836), .B(n844), .Y(n832) );
  NAND2X1 U490 ( .A(n1050), .B(n1123), .Y(n837) );
  AND2X2 U491 ( .A(n1074), .B(n849), .Y(n692) );
  NAND2X2 U492 ( .A(counterRead[1]), .B(n1092), .Y(n828) );
  INVX3 U493 ( .A(n840), .Y(n818) );
  NAND2X1 U494 ( .A(n801), .B(n849), .Y(n807) );
  CLKINVX1 U495 ( .A(n804), .Y(n813) );
  NAND2X1 U496 ( .A(n700), .B(n746), .Y(n849) );
  CLKAND2X3 U497 ( .A(n101), .B(n494), .Y(n700) );
  NAND2X1 U498 ( .A(counterRead[1]), .B(n494), .Y(n804) );
  CLKINVX1 U499 ( .A(counterRead[1]), .Y(n746) );
  NAND2X6 U500 ( .A(n101), .B(n818), .Y(n1072) );
  NAND2X2 U501 ( .A(n684), .B(n1006), .Y(n844) );
  NAND2X1 U502 ( .A(n813), .B(n101), .Y(n845) );
  NAND2X1 U503 ( .A(n813), .B(n719), .Y(n801) );
  NAND2BX1 U504 ( .AN(N610), .B(n1079), .Y(n1010) );
  INVX16 U505 ( .A(n707), .Y(n1123) );
  NAND3BX1 U506 ( .AN(n78), .B(n471), .C(n759), .Y(n1054) );
  BUFX4 U507 ( .A(mulTemp[15]), .Y(n558) );
  INVX3 U508 ( .A(n99), .Y(n1006) );
  BUFX8 U509 ( .A(counterRead[0]), .Y(n719) );
  CLKBUFX3 U510 ( .A(mulTemp[6]), .Y(n557) );
  NAND2X1 U511 ( .A(n1093), .B(n1095), .Y(n1094) );
  NAND3BX1 U512 ( .AN(n1023), .B(n1016), .C(n1015), .Y(n371) );
  CLKINVX1 U513 ( .A(mulTemp[30]), .Y(n874) );
  AOI2BB2X1 U514 ( .B0(N735), .B1(n1036), .A0N(n720), .A1N(n866), .Y(n869) );
  AND2X2 U515 ( .A(n1066), .B(n1052), .Y(n472) );
  AOI21X2 U516 ( .A0(n294), .A1(n784), .B0(n786), .Y(n473) );
  AO22X1 U517 ( .A0(n1135), .A1(n1108), .B0(n716), .B1(n142), .Y(n474) );
  OR3X2 U518 ( .A(n502), .B(n503), .C(n504), .Y(n475) );
  OR3X2 U519 ( .A(n505), .B(n506), .C(n507), .Y(n476) );
  OR3X2 U520 ( .A(n508), .B(n509), .C(n510), .Y(n477) );
  OR3X2 U521 ( .A(n511), .B(n512), .C(n513), .Y(n478) );
  OR3X2 U522 ( .A(n514), .B(n515), .C(n516), .Y(n479) );
  OR3X2 U523 ( .A(n517), .B(n518), .C(n519), .Y(n480) );
  OR3X2 U524 ( .A(n520), .B(n521), .C(n522), .Y(n481) );
  OR3X2 U525 ( .A(n523), .B(n524), .C(n525), .Y(n482) );
  OR3X2 U526 ( .A(n526), .B(n527), .C(n528), .Y(n483) );
  OR3X2 U527 ( .A(n529), .B(n530), .C(n531), .Y(n484) );
  OR3X2 U528 ( .A(n532), .B(n533), .C(n534), .Y(n485) );
  OR3X2 U529 ( .A(n535), .B(n536), .C(n537), .Y(n486) );
  OR3X2 U530 ( .A(n538), .B(n539), .C(n540), .Y(n487) );
  OR3X2 U531 ( .A(n541), .B(n542), .C(n543), .Y(n488) );
  OR3X2 U532 ( .A(n544), .B(n545), .C(n546), .Y(n489) );
  OR3X2 U533 ( .A(n547), .B(n548), .C(n549), .Y(n490) );
  OR3X2 U534 ( .A(n550), .B(n551), .C(n552), .Y(n491) );
  OR3X2 U535 ( .A(n553), .B(n554), .C(n555), .Y(n492) );
  AND3X2 U536 ( .A(n845), .B(n844), .C(n814), .Y(n493) );
  OAI211X1 U537 ( .A0(n798), .A1(n797), .B0(n811), .C0(n840), .Y(n816) );
  AND2X4 U538 ( .A(n743), .B(n805), .Y(n494) );
  CLKAND2X3 U539 ( .A(n706), .B(n742), .Y(n495) );
  AOI21X1 U540 ( .A0(n693), .A1(n694), .B0(n760), .Y(n496) );
  OR4X1 U541 ( .A(n192), .B(n712), .C(n716), .D(n715), .Y(n497) );
  INVX3 U542 ( .A(n846), .Y(n1092) );
  INVX4 U543 ( .A(counterRead[3]), .Y(n805) );
  INVX12 U544 ( .A(n498), .Y(cwr) );
  INVX12 U546 ( .A(n500), .Y(crd) );
  CLKINVX1 U547 ( .A(n138), .Y(n1122) );
  AND2X2 U548 ( .A(n1137), .B(n709), .Y(n502) );
  AND2XL U549 ( .A(cdata_rd[18]), .B(n710), .Y(n503) );
  AND2X2 U550 ( .A(roundTemp[19]), .B(n711), .Y(n504) );
  AND2X2 U551 ( .A(n1138), .B(n709), .Y(n505) );
  AND2XL U552 ( .A(cdata_rd[17]), .B(n710), .Y(n506) );
  AND2X2 U553 ( .A(roundTemp[18]), .B(n711), .Y(n507) );
  AND2X2 U554 ( .A(n1139), .B(n709), .Y(n508) );
  AND2XL U555 ( .A(cdata_rd[16]), .B(n710), .Y(n509) );
  AND2X2 U556 ( .A(roundTemp[17]), .B(n711), .Y(n510) );
  AND2X2 U557 ( .A(n1140), .B(n709), .Y(n511) );
  AND2XL U558 ( .A(cdata_rd[15]), .B(n710), .Y(n512) );
  AND2X2 U559 ( .A(roundTemp[16]), .B(n711), .Y(n513) );
  AND2X2 U560 ( .A(n1141), .B(n709), .Y(n514) );
  AND2XL U561 ( .A(cdata_rd[14]), .B(n710), .Y(n515) );
  AND2X2 U562 ( .A(roundTemp[15]), .B(n711), .Y(n516) );
  AND2X2 U563 ( .A(n1142), .B(n709), .Y(n517) );
  AND2XL U564 ( .A(cdata_rd[13]), .B(n710), .Y(n518) );
  AND2X2 U565 ( .A(roundTemp[14]), .B(n711), .Y(n519) );
  AND2X2 U566 ( .A(n1143), .B(n709), .Y(n520) );
  AND2XL U567 ( .A(cdata_rd[12]), .B(n710), .Y(n521) );
  AND2X2 U568 ( .A(roundTemp[13]), .B(n711), .Y(n522) );
  AND2X2 U569 ( .A(n1144), .B(n709), .Y(n523) );
  AND2XL U570 ( .A(cdata_rd[11]), .B(n710), .Y(n524) );
  AND2X2 U571 ( .A(roundTemp[12]), .B(n711), .Y(n525) );
  AND2X2 U572 ( .A(n1145), .B(n709), .Y(n526) );
  AND2XL U573 ( .A(cdata_rd[10]), .B(n710), .Y(n527) );
  AND2X2 U574 ( .A(roundTemp[11]), .B(n711), .Y(n528) );
  AND2X2 U575 ( .A(n1146), .B(n709), .Y(n529) );
  AND2XL U576 ( .A(cdata_rd[9]), .B(n710), .Y(n530) );
  AND2X2 U577 ( .A(roundTemp[10]), .B(n711), .Y(n531) );
  AND2X2 U578 ( .A(n1147), .B(n709), .Y(n532) );
  AND2XL U579 ( .A(cdata_rd[8]), .B(n710), .Y(n533) );
  AND2X2 U580 ( .A(roundTemp[9]), .B(n711), .Y(n534) );
  AND2X2 U581 ( .A(n1148), .B(n709), .Y(n535) );
  AND2XL U582 ( .A(cdata_rd[7]), .B(n710), .Y(n536) );
  AND2X2 U583 ( .A(roundTemp[8]), .B(n711), .Y(n537) );
  AND2X2 U584 ( .A(n1149), .B(n709), .Y(n538) );
  AND2XL U585 ( .A(cdata_rd[6]), .B(n710), .Y(n539) );
  AND2X2 U586 ( .A(roundTemp[7]), .B(n711), .Y(n540) );
  AND2X2 U587 ( .A(n1150), .B(n709), .Y(n541) );
  AND2XL U588 ( .A(cdata_rd[5]), .B(n710), .Y(n542) );
  AND2X2 U589 ( .A(roundTemp[6]), .B(n711), .Y(n543) );
  AND2X2 U590 ( .A(n1151), .B(n709), .Y(n544) );
  AND2XL U591 ( .A(cdata_rd[4]), .B(n710), .Y(n545) );
  AND2X2 U592 ( .A(roundTemp[5]), .B(n711), .Y(n546) );
  AND2X2 U593 ( .A(n1152), .B(n709), .Y(n547) );
  AND2XL U594 ( .A(cdata_rd[3]), .B(n710), .Y(n548) );
  AND2X2 U595 ( .A(roundTemp[4]), .B(n711), .Y(n549) );
  AND2X2 U596 ( .A(n1153), .B(n709), .Y(n550) );
  AND2XL U597 ( .A(cdata_rd[2]), .B(n710), .Y(n551) );
  AND2X2 U598 ( .A(roundTemp[3]), .B(n711), .Y(n552) );
  AND2X2 U599 ( .A(n1154), .B(n709), .Y(n553) );
  AND2XL U600 ( .A(cdata_rd[1]), .B(n710), .Y(n554) );
  AND2X2 U601 ( .A(roundTemp[2]), .B(n711), .Y(n555) );
  OA21X4 U602 ( .A0(n1123), .A1(n825), .B0(n843), .Y(n556) );
  NAND2X4 U603 ( .A(n556), .B(n845), .Y(kernelTemp[5]) );
  INVXL U604 ( .A(n832), .Y(n825) );
  NAND2X6 U605 ( .A(n818), .B(n719), .Y(n843) );
  NAND2X2 U606 ( .A(n493), .B(n687), .Y(kernelTemp[10]) );
  NAND4BX2 U607 ( .AN(n817), .B(n833), .C(n812), .D(n814), .Y(kernelTemp[11])
         );
  NAND3X2 U608 ( .A(n814), .B(n796), .C(n830), .Y(kernelTemp[19]) );
  INVX2 U609 ( .A(n98), .Y(n743) );
  NAND2X2 U610 ( .A(n837), .B(n800), .Y(kernelTemp[15]) );
  MXI2X1 U611 ( .A(n799), .B(n816), .S0(n1123), .Y(n800) );
  BUFX4 U612 ( .A(n826), .Y(n559) );
  NAND2XL U613 ( .A(n99), .B(n494), .Y(n826) );
  MXI2X1 U614 ( .A(n799), .B(n818), .S0(n1123), .Y(n796) );
  OAI21X1 U615 ( .A0(n832), .A1(n831), .B0(n707), .Y(n834) );
  BUFX6 U616 ( .A(mulTemp[28]), .Y(n560) );
  BUFX6 U617 ( .A(n1100), .Y(n561) );
  NAND2XL U618 ( .A(n1072), .B(n804), .Y(n1100) );
  OAI211X4 U619 ( .A0(n819), .A1(n1123), .B0(n837), .C0(n1072), .Y(
        kernelTemp[7]) );
  INVXL U620 ( .A(mulTemp[17]), .Y(n926) );
  NAND2X2 U621 ( .A(n101), .B(n699), .Y(n811) );
  NAND2X8 U622 ( .A(n719), .B(n1050), .Y(n1076) );
  NAND2XL U623 ( .A(n719), .B(n494), .Y(n836) );
  NAND2X2 U624 ( .A(n684), .B(n1123), .Y(n830) );
  AND2X1 U625 ( .A(n101), .B(n699), .Y(n684) );
  INVX12 U626 ( .A(n562), .Y(cdata_wr[16]) );
  INVX12 U627 ( .A(n564), .Y(cdata_wr[7]) );
  INVX12 U628 ( .A(n566), .Y(cdata_wr[1]) );
  INVX12 U629 ( .A(n568), .Y(cdata_wr[2]) );
  INVX12 U630 ( .A(n570), .Y(cdata_wr[10]) );
  INVX12 U631 ( .A(n572), .Y(cdata_wr[14]) );
  INVX12 U632 ( .A(n574), .Y(cdata_wr[17]) );
  OAI211XL U633 ( .A0(n81), .A1(n1067), .B0(n1066), .C0(n1065), .Y(N430) );
  BUFX12 U634 ( .A(n1133), .Y(iaddr[6]) );
  INVX12 U635 ( .A(n578), .Y(iaddr[0]) );
  INVX12 U636 ( .A(n580), .Y(busy) );
  INVX12 U637 ( .A(n582), .Y(iaddr[8]) );
  INVX12 U639 ( .A(n586), .Y(iaddr[2]) );
  INVX12 U640 ( .A(n588), .Y(iaddr[1]) );
  INVX12 U641 ( .A(n590), .Y(caddr_rd[9]) );
  INVX12 U642 ( .A(n592), .Y(caddr_rd[8]) );
  INVX12 U643 ( .A(n594), .Y(caddr_rd[7]) );
  INVX12 U644 ( .A(n596), .Y(caddr_rd[6]) );
  INVX12 U645 ( .A(n598), .Y(caddr_rd[5]) );
  INVX12 U646 ( .A(n600), .Y(caddr_rd[4]) );
  INVX12 U647 ( .A(n602), .Y(caddr_rd[3]) );
  INVX12 U648 ( .A(n604), .Y(caddr_rd[2]) );
  INVX12 U649 ( .A(n606), .Y(caddr_rd[1]) );
  INVX12 U650 ( .A(n608), .Y(caddr_rd[0]) );
  INVX12 U651 ( .A(n610), .Y(caddr_wr[10]) );
  INVX12 U652 ( .A(n612), .Y(caddr_wr[5]) );
  INVX12 U653 ( .A(n614), .Y(caddr_wr[4]) );
  INVX12 U654 ( .A(n616), .Y(caddr_wr[3]) );
  INVX12 U655 ( .A(n618), .Y(caddr_wr[2]) );
  INVX12 U656 ( .A(n620), .Y(caddr_wr[1]) );
  INVX12 U657 ( .A(n622), .Y(iaddr[9]) );
  INVX12 U658 ( .A(n624), .Y(iaddr[3]) );
  INVX12 U659 ( .A(n626), .Y(caddr_wr[9]) );
  INVX12 U660 ( .A(n628), .Y(caddr_wr[8]) );
  INVX12 U661 ( .A(n630), .Y(caddr_wr[7]) );
  INVX12 U662 ( .A(n632), .Y(caddr_wr[6]) );
  INVX12 U663 ( .A(n634), .Y(iaddr[11]) );
  INVX12 U664 ( .A(n636), .Y(iaddr[10]) );
  INVX12 U665 ( .A(n638), .Y(iaddr[5]) );
  INVX12 U666 ( .A(n640), .Y(iaddr[4]) );
  INVX12 U667 ( .A(n642), .Y(caddr_wr[0]) );
  INVX12 U668 ( .A(n644), .Y(caddr_rd[11]) );
  INVX12 U669 ( .A(n646), .Y(caddr_rd[10]) );
  INVX12 U670 ( .A(n648), .Y(csel[1]) );
  INVX12 U671 ( .A(n650), .Y(csel[2]) );
  INVX12 U672 ( .A(n652), .Y(csel[0]) );
  INVX12 U673 ( .A(n654), .Y(caddr_wr[11]) );
  INVX12 U674 ( .A(n656), .Y(cdata_wr[15]) );
  INVX12 U675 ( .A(n658), .Y(cdata_wr[6]) );
  INVX12 U676 ( .A(n660), .Y(cdata_wr[13]) );
  INVX12 U677 ( .A(n662), .Y(cdata_wr[11]) );
  INVX12 U678 ( .A(n664), .Y(cdata_wr[4]) );
  INVX12 U679 ( .A(n666), .Y(cdata_wr[9]) );
  INVX12 U680 ( .A(n668), .Y(cdata_wr[0]) );
  INVX12 U681 ( .A(n670), .Y(cdata_wr[18]) );
  INVX12 U682 ( .A(n672), .Y(cdata_wr[3]) );
  INVX12 U683 ( .A(n674), .Y(cdata_wr[8]) );
  INVX12 U684 ( .A(n676), .Y(cdata_wr[5]) );
  INVX12 U685 ( .A(n678), .Y(cdata_wr[19]) );
  INVX12 U686 ( .A(n680), .Y(cdata_wr[12]) );
  INVX12 U687 ( .A(n828), .Y(n1050) );
  NAND2X6 U688 ( .A(n699), .B(n99), .Y(n840) );
  AND2XL U689 ( .A(n700), .B(n746), .Y(n682) );
  NAND2X2 U690 ( .A(n92), .B(n98), .Y(n846) );
  NAND2BX2 U691 ( .AN(n559), .B(n719), .Y(n1073) );
  INVXL U692 ( .A(n1092), .Y(n683) );
  NAND3BX4 U693 ( .AN(n838), .B(n691), .C(n837), .Y(kernelTemp[2]) );
  AND2XL U694 ( .A(n471), .B(current_State[3]), .Y(n705) );
  AND2X1 U695 ( .A(n836), .B(n1074), .Y(n691) );
  CLKINVX2 U696 ( .A(n92), .Y(n798) );
  NAND2X6 U697 ( .A(n719), .B(counterRead[1]), .Y(n1091) );
  NAND2X1 U698 ( .A(n101), .B(counterRead[1]), .Y(n797) );
  NAND2XL U699 ( .A(n700), .B(n1123), .Y(n823) );
  INVXL U700 ( .A(mulTemp[26]), .Y(n890) );
  NAND2XL U701 ( .A(n820), .B(n1072), .Y(n821) );
  AND2X1 U702 ( .A(n809), .B(n840), .Y(n690) );
  BUFX20 U703 ( .A(BiasTemp_7), .Y(n707) );
  NOR2BX4 U704 ( .AN(n798), .B(counterRead[2]), .Y(n699) );
  INVX1 U705 ( .A(mulTemp[16]), .Y(n930) );
  INVX1 U706 ( .A(mulTemp[29]), .Y(n878) );
  INVX1 U707 ( .A(n560), .Y(n882) );
  INVX1 U708 ( .A(mulTemp[27]), .Y(n886) );
  INVXL U709 ( .A(n558), .Y(n934) );
  INVXL U710 ( .A(mulTemp[9]), .Y(n958) );
  INVXL U711 ( .A(mulTemp[13]), .Y(n942) );
  CLKINVX1 U712 ( .A(mulTemp[8]), .Y(n962) );
  INVXL U713 ( .A(mulTemp[5]), .Y(n974) );
  INVX1 U714 ( .A(mulTemp[12]), .Y(n946) );
  INVX1 U715 ( .A(mulTemp[11]), .Y(n950) );
  NAND2X6 U716 ( .A(n685), .B(n80), .Y(BiasTemp_7) );
  NAND4XL U717 ( .A(n835), .B(n830), .C(n829), .D(n828), .Y(kernelTemp[4]) );
  AOI2BB2X1 U718 ( .B0(N734), .B1(n724), .A0N(n720), .A1N(n870), .Y(n873) );
  AOI2BB2X1 U719 ( .B0(N740), .B1(n724), .A0N(n1031), .A1N(n1027), .Y(n1030)
         );
  AOI2BB2X1 U720 ( .B0(N741), .B1(n724), .A0N(n721), .A1N(n1027), .Y(n1026) );
  AOI2BB2X1 U721 ( .B0(N737), .B1(n724), .A0N(n720), .A1N(n998), .Y(n1001) );
  AOI2BB2X1 U722 ( .B0(N738), .B1(n724), .A0N(n721), .A1N(n1002), .Y(n1005) );
  AOI2BB2X1 U723 ( .B0(N736), .B1(n725), .A0N(n720), .A1N(n861), .Y(n865) );
  AOI2BB2X1 U724 ( .B0(N727), .B1(n726), .A0N(n720), .A1N(n898), .Y(n901) );
  NAND2X1 U725 ( .A(N744), .B(n1036), .Y(n1016) );
  NAND2X1 U726 ( .A(N743), .B(n726), .Y(n1019) );
  NAND2X1 U727 ( .A(N745), .B(n725), .Y(n1013) );
  AOI2BB2X1 U728 ( .B0(N725), .B1(n726), .A0N(n720), .A1N(n906), .Y(n909) );
  AOI2BB2X1 U729 ( .B0(N724), .B1(n726), .A0N(n721), .A1N(n910), .Y(n913) );
  AOI2BB2X1 U730 ( .B0(N726), .B1(n726), .A0N(n720), .A1N(n902), .Y(n905) );
  INVXL U731 ( .A(n685), .Y(n853) );
  INVX1 U732 ( .A(current_State[0]), .Y(n759) );
  INVXL U733 ( .A(mulTemp[21]), .Y(n910) );
  INVXL U734 ( .A(mulTemp[34]), .Y(n998) );
  INVXL U735 ( .A(mulTemp[31]), .Y(n870) );
  INVXL U736 ( .A(mulTemp[18]), .Y(n922) );
  INVXL U737 ( .A(mulTemp[19]), .Y(n918) );
  INVXL U738 ( .A(mulTemp[25]), .Y(n894) );
  INVXL U739 ( .A(mulTemp[10]), .Y(n954) );
  INVXL U740 ( .A(mulTemp[7]), .Y(n966) );
  INVXL U741 ( .A(mulTemp[2]), .Y(n986) );
  INVX1 U742 ( .A(n557), .Y(n970) );
  INVXL U743 ( .A(mulTemp[4]), .Y(n978) );
  MX2XL U744 ( .A(n690), .B(n1076), .S0(n1123), .Y(n810) );
  INVXL U745 ( .A(n801), .Y(n851) );
  CLKINVX1 U746 ( .A(n1037), .Y(n1033) );
  NAND2XL U747 ( .A(n806), .B(n699), .Y(n771) );
  CLKINVX1 U748 ( .A(n859), .Y(n1036) );
  NAND2XL U749 ( .A(n844), .B(n845), .Y(n856) );
  NAND4XL U750 ( .A(n1080), .B(n1076), .C(n843), .D(n1072), .Y(n858) );
  INVXL U751 ( .A(n1074), .Y(n860) );
  NAND3BXL U752 ( .AN(n1006), .B(n719), .C(n1092), .Y(n1079) );
  NAND3BXL U753 ( .AN(counterRead[3]), .B(n1123), .C(n1006), .Y(n829) );
  NAND3BX2 U754 ( .AN(n1040), .B(n1039), .C(n1038), .Y(n369) );
  AO22X4 U755 ( .A0(N1107), .A1(n728), .B0(N746), .B1(n725), .Y(n1040) );
  AOI32XL U756 ( .A0(ready), .A1(n78), .A2(n759), .B0(n771), .B1(n1123), .Y(
        n766) );
  AOI32XL U757 ( .A0(current_State[0]), .A1(current_State[3]), .A2(n704), .B0(
        n682), .B1(n770), .Y(n774) );
  OA22XL U758 ( .A0(n707), .A1(n771), .B0(n776), .B1(n1070), .Y(n773) );
  OAI31XL U759 ( .A0(n719), .A1(counterRead[1]), .A2(n683), .B0(n845), .Y(
        n1075) );
  NAND2X2 U760 ( .A(n1009), .B(current_State[1]), .Y(n1071) );
  NAND2XL U761 ( .A(n80), .B(current_State[0]), .Y(n744) );
  AND2XL U762 ( .A(current_State[1]), .B(current_State[0]), .Y(n701) );
  OAI32XL U763 ( .A0(counterRead[2]), .A1(n1091), .A2(n757), .B0(n98), .B1(
        n756), .Y(n465) );
  MXI2XL U764 ( .A(n1094), .B(n1101), .S0(N314), .Y(n703) );
  NAND2XL U765 ( .A(n80), .B(n471), .Y(n1067) );
  CLKINVX1 U766 ( .A(mulTemp[24]), .Y(n898) );
  CLKINVX1 U767 ( .A(mulTemp[23]), .Y(n902) );
  CLKINVX1 U768 ( .A(mulTemp[22]), .Y(n906) );
  CLKINVX1 U769 ( .A(mulTemp[35]), .Y(n1002) );
  CLKINVX1 U770 ( .A(mulTemp[32]), .Y(n866) );
  CLKINVX1 U771 ( .A(mulTemp[37]), .Y(n1027) );
  CLKINVX1 U772 ( .A(mulTemp[20]), .Y(n914) );
  CLKINVX1 U773 ( .A(mulTemp[14]), .Y(n938) );
  CLKINVX1 U774 ( .A(mulTemp[3]), .Y(n982) );
  CLKBUFX3 U775 ( .A(n686), .Y(n727) );
  CLKBUFX3 U776 ( .A(n686), .Y(n728) );
  CLKINVX1 U777 ( .A(n807), .Y(n1080) );
  INVX3 U778 ( .A(n793), .Y(n1109) );
  AND2X2 U779 ( .A(n722), .B(n862), .Y(n686) );
  CLKBUFX3 U780 ( .A(n1033), .Y(n722) );
  CLKINVX1 U781 ( .A(mulTemp[1]), .Y(n990) );
  NAND2X1 U782 ( .A(n1111), .B(n786), .Y(n277) );
  NOR2BX2 U783 ( .AN(n285), .B(n1111), .Y(n287) );
  NAND2X1 U784 ( .A(n752), .B(n751), .Y(n748) );
  CLKINVX1 U785 ( .A(n789), .Y(n770) );
  CLKBUFX3 U786 ( .A(n1033), .Y(n723) );
  CLKINVX1 U787 ( .A(mulTemp[0]), .Y(n994) );
  CLKBUFX3 U788 ( .A(n1031), .Y(n720) );
  CLKBUFX3 U789 ( .A(n1031), .Y(n721) );
  CLKINVX1 U790 ( .A(n1060), .Y(n1106) );
  CLKBUFX3 U791 ( .A(n731), .Y(n736) );
  CLKBUFX3 U792 ( .A(n731), .Y(n733) );
  CLKBUFX3 U793 ( .A(n731), .Y(n734) );
  CLKBUFX3 U794 ( .A(n731), .Y(n737) );
  CLKBUFX3 U795 ( .A(n731), .Y(n735) );
  CLKBUFX3 U796 ( .A(n731), .Y(n738) );
  CLKBUFX3 U797 ( .A(n731), .Y(n741) );
  CLKBUFX3 U798 ( .A(n731), .Y(n739) );
  CLKBUFX3 U799 ( .A(n731), .Y(n740) );
  CLKBUFX3 U800 ( .A(n731), .Y(n732) );
  CLKINVX1 U801 ( .A(n835), .Y(n838) );
  NAND2X1 U802 ( .A(n1073), .B(n810), .Y(kernelTemp[12]) );
  NAND3X1 U803 ( .A(n833), .B(n808), .C(n830), .Y(kernelTemp[13]) );
  MXI2X1 U804 ( .A(n815), .B(n807), .S0(n1123), .Y(n808) );
  CLKINVX1 U805 ( .A(n561), .Y(n1093) );
  NAND2X1 U806 ( .A(n824), .B(n823), .Y(kernelTemp[6]) );
  MXI2X1 U807 ( .A(n822), .B(n821), .S0(n1123), .Y(n824) );
  NAND2X1 U808 ( .A(n690), .B(n1073), .Y(n822) );
  NAND2X1 U809 ( .A(n790), .B(n1053), .Y(n793) );
  AND4X1 U810 ( .A(n698), .B(n1109), .C(n472), .D(n696), .Y(n264) );
  CLKINVX1 U811 ( .A(n1039), .Y(n1023) );
  CLKBUFX3 U812 ( .A(n729), .Y(n742) );
  CLKBUFX3 U813 ( .A(n730), .Y(n729) );
  INVX3 U814 ( .A(n142), .Y(n1111) );
  CLKINVX1 U815 ( .A(n780), .Y(n1110) );
  CLKINVX1 U816 ( .A(n771), .Y(n862) );
  CLKBUFX3 U817 ( .A(n1036), .Y(n726) );
  CLKBUFX3 U818 ( .A(n1036), .Y(n725) );
  CLKBUFX3 U819 ( .A(n1036), .Y(n724) );
  AND2X2 U820 ( .A(n769), .B(n1052), .Y(n775) );
  NOR2X2 U821 ( .A(n1111), .B(n1113), .Y(n279) );
  OAI2BB1X1 U822 ( .A0N(n785), .A1N(n783), .B0(n784), .Y(n285) );
  NAND2X1 U823 ( .A(n768), .B(n693), .Y(n789) );
  NAND2X1 U824 ( .A(n142), .B(n1113), .Y(n784) );
  NAND2X1 U825 ( .A(n688), .B(n757), .Y(n751) );
  NAND2X1 U826 ( .A(n750), .B(n101), .Y(n752) );
  NAND2BX1 U827 ( .AN(n748), .B(n749), .Y(n755) );
  CLKINVX1 U828 ( .A(n1087), .Y(n1078) );
  CLKINVX1 U829 ( .A(n1073), .Y(n857) );
  CLKINVX1 U830 ( .A(n757), .Y(n750) );
  CLKINVX1 U831 ( .A(n781), .Y(n764) );
  AOI21X1 U832 ( .A0(n682), .A1(n1049), .B0(n862), .Y(n688) );
  CLKINVX1 U833 ( .A(n1105), .Y(n760) );
  CLKINVX1 U834 ( .A(n351), .Y(n1124) );
  NAND2X1 U835 ( .A(n1050), .B(n1049), .Y(n1063) );
  NAND2X1 U836 ( .A(n1080), .B(n1079), .Y(n1088) );
  NAND2X2 U837 ( .A(n1007), .B(n472), .Y(n1060) );
  CLKINVX1 U838 ( .A(n1049), .Y(n1007) );
  AND2X2 U839 ( .A(n1092), .B(n1049), .Y(n689) );
  CLKINVX1 U840 ( .A(n785), .Y(n786) );
  CLKINVX1 U841 ( .A(n1095), .Y(n1102) );
  AO21X1 U842 ( .A0(n1010), .A1(n1049), .B0(n1009), .Y(n118) );
  MXI2X1 U843 ( .A(n1010), .B(n1008), .S0(n1007), .Y(n117) );
  NAND2X1 U844 ( .A(n1054), .B(n1111), .Y(n1008) );
  NAND2BX1 U845 ( .AN(n809), .B(n1123), .Y(n833) );
  CLKINVX1 U846 ( .A(n1101), .Y(n819) );
  NAND2X1 U847 ( .A(n1072), .B(n839), .Y(kernelTemp[1]) );
  CLKMX2X2 U848 ( .A(n1076), .B(n692), .S0(n1123), .Y(n839) );
  CLKMX2X2 U849 ( .A(n811), .B(n843), .S0(n1123), .Y(n812) );
  NAND2X1 U850 ( .A(n843), .B(n803), .Y(kernelTemp[14]) );
  CLKMX2X2 U851 ( .A(n802), .B(n1080), .S0(n1123), .Y(n803) );
  AND2X2 U852 ( .A(n809), .B(n559), .Y(n802) );
  CLKMX2X2 U853 ( .A(n816), .B(n815), .S0(n1123), .Y(kernelTemp[9]) );
  CLKMX2X2 U854 ( .A(n827), .B(n840), .S0(n1123), .Y(n835) );
  AND2X2 U855 ( .A(n1072), .B(n559), .Y(n827) );
  NAND2X1 U856 ( .A(n687), .B(n842), .Y(kernelTemp[0]) );
  CLKMX2X2 U857 ( .A(n841), .B(n1076), .S0(n1123), .Y(n842) );
  AND2X2 U858 ( .A(n691), .B(n840), .Y(n841) );
  CLKBUFX3 U859 ( .A(n1103), .Y(n706) );
  CLKINVX1 U860 ( .A(n853), .Y(n1103) );
  NAND2X1 U861 ( .A(n834), .B(n833), .Y(kernelTemp[3]) );
  CLKINVX1 U862 ( .A(n843), .Y(n831) );
  AO21X1 U863 ( .A0(n818), .A1(n707), .B0(n817), .Y(kernelTemp[8]) );
  NAND4X1 U864 ( .A(next_State[0]), .B(n779), .C(next_State[1]), .D(
        next_State[2]), .Y(n790) );
  CLKINVX1 U865 ( .A(next_State[3]), .Y(n779) );
  NAND4BBXL U866 ( .AN(next_State[0]), .BN(next_State[2]), .C(next_State[3]), 
        .D(next_State[1]), .Y(n1053) );
  NAND3BX1 U867 ( .AN(n1074), .B(mulTemp_43), .C(n722), .Y(n1039) );
  CLKINVX1 U868 ( .A(n1091), .Y(n806) );
  NAND2X1 U869 ( .A(n209), .B(n210), .Y(n421) );
  AOI222XL U870 ( .A0(n712), .A1(n793), .B0(n714), .B1(n142), .C0(n792), .C1(
        n713), .Y(n210) );
  OA22X1 U871 ( .A0(n708), .A1(n630), .B0(n45), .B1(n1071), .Y(n209) );
  NAND2X1 U872 ( .A(n211), .B(n212), .Y(n422) );
  AOI222XL U873 ( .A0(n792), .A1(n712), .B0(n715), .B1(n793), .C0(n713), .C1(
        n142), .Y(n212) );
  OA22X1 U874 ( .A0(n708), .A1(n628), .B0(n44), .B1(n1071), .Y(n211) );
  NAND2X1 U875 ( .A(n213), .B(n214), .Y(n423) );
  AOI222XL U876 ( .A0(n712), .A1(n142), .B0(n716), .B1(n793), .C0(n792), .C1(
        n715), .Y(n214) );
  OA22X1 U877 ( .A0(n708), .A1(n626), .B0(n43), .B1(n1071), .Y(n213) );
  CLKBUFX3 U878 ( .A(n1068), .Y(n708) );
  NAND3BX1 U879 ( .AN(n780), .B(n1109), .C(n1071), .Y(n1068) );
  NAND2X1 U880 ( .A(n790), .B(n1066), .Y(n1051) );
  NAND3BX1 U881 ( .AN(n142), .B(n1109), .C(n1054), .Y(N422) );
  CLKBUFX3 U882 ( .A(n1112), .Y(n730) );
  NAND2X1 U883 ( .A(n1070), .B(n1111), .Y(n780) );
  AND2X2 U884 ( .A(n759), .B(current_State[1]), .Y(n694) );
  OAI221XL U885 ( .A0(n1072), .A1(n850), .B0(n1113), .B1(n844), .C0(n843), .Y(
        n848) );
  OAI211X1 U886 ( .A0(n351), .A1(n787), .B0(n778), .C0(n777), .Y(next_State[2]) );
  AND4X1 U887 ( .A(n695), .B(n496), .C(n472), .D(n789), .Y(n777) );
  AOI32X1 U888 ( .A0(n862), .A1(n706), .A2(current_State[1]), .B0(n776), .B1(
        n792), .Y(n778) );
  OAI31XL U889 ( .A0(n858), .A1(n857), .A2(n856), .B0(n722), .Y(n859) );
  CLKINVX1 U890 ( .A(n1054), .Y(n1009) );
  CLKINVX1 U891 ( .A(n1070), .Y(n792) );
  AO21X1 U892 ( .A0(n855), .A1(n854), .B0(n853), .Y(n1037) );
  AOI222XL U893 ( .A0(n857), .A1(n184), .B0(n852), .B1(n497), .C0(n851), .C1(
        n191), .Y(n854) );
  AOI211X1 U894 ( .A0(n848), .A1(n847), .B0(n862), .C0(n1075), .Y(n855) );
  CLKINVX1 U895 ( .A(n1071), .Y(n795) );
  CLKINVX1 U896 ( .A(n762), .Y(n769) );
  OAI211X1 U897 ( .A0(n782), .A1(n763), .B0(n496), .C0(n761), .Y(n762) );
  NAND3BX1 U898 ( .AN(n862), .B(n706), .C(current_State[1]), .Y(n761) );
  CLKINVX1 U899 ( .A(n294), .Y(n783) );
  AOI21X1 U900 ( .A0(n764), .A1(n763), .B0(n795), .Y(n695) );
  NAND3X1 U901 ( .A(n1072), .B(n1074), .C(n1073), .Y(n1087) );
  NAND2X1 U902 ( .A(n1065), .B(n789), .Y(n1049) );
  NAND3BX1 U903 ( .AN(n1009), .B(n782), .C(n781), .Y(n785) );
  OAI221XL U904 ( .A0(n850), .A1(n1074), .B0(n1113), .B1(n849), .C0(n1076), 
        .Y(n852) );
  NAND2X1 U905 ( .A(n722), .B(n860), .Y(n1031) );
  NAND2X1 U906 ( .A(n688), .B(n745), .Y(n757) );
  NAND2X1 U907 ( .A(n768), .B(n705), .Y(n1052) );
  CLKINVX1 U908 ( .A(n191), .Y(n1113) );
  NAND2X1 U909 ( .A(n693), .B(n701), .Y(n781) );
  NAND2X1 U910 ( .A(n750), .B(n746), .Y(n749) );
  NAND2X1 U911 ( .A(n705), .B(n701), .Y(n1105) );
  NAND2X1 U912 ( .A(n1113), .B(n185), .Y(n351) );
  CLKINVX1 U913 ( .A(n763), .Y(n776) );
  CLKINVX1 U914 ( .A(n1065), .Y(n758) );
  NAND2BX1 U915 ( .AN(n1075), .B(n1076), .Y(n1089) );
  CLKINVX1 U916 ( .A(n184), .Y(n850) );
  CLKINVX1 U917 ( .A(n744), .Y(n768) );
  AO22X1 U918 ( .A0(n747), .A1(n719), .B0(n748), .B1(n1006), .Y(n466) );
  CLKINVX1 U919 ( .A(n749), .Y(n747) );
  AO22X1 U920 ( .A0(n750), .A1(n851), .B0(n755), .B1(n798), .Y(n467) );
  CLKINVX1 U921 ( .A(n185), .Y(n847) );
  NAND2X1 U922 ( .A(n689), .B(n719), .Y(n1048) );
  AND3X2 U923 ( .A(n788), .B(n789), .C(n1054), .Y(n696) );
  AND2X2 U924 ( .A(n294), .B(n785), .Y(n697) );
  AND2X2 U925 ( .A(n1065), .B(n787), .Y(n698) );
  ADDHX1 U926 ( .A(n713), .B(\r363/carry[2] ), .CO(\r363/carry[3] ), .S(
        index_Y_After[2]) );
  ADDHX1 U927 ( .A(n712), .B(\r363/carry[3] ), .CO(\r363/carry[4] ), .S(
        index_Y_After[3]) );
  ADDHX1 U928 ( .A(n717), .B(\r361/carry[3] ), .CO(\r361/carry[4] ), .S(
        index_X_After[3]) );
  AO21X1 U929 ( .A0(n754), .A1(n719), .B0(n753), .Y(n468) );
  CLKINVX1 U930 ( .A(n751), .Y(n754) );
  CLKINVX1 U931 ( .A(n752), .Y(n753) );
  ADDHX1 U932 ( .A(n715), .B(\r363/carry[4] ), .CO(\r363/carry[5] ), .S(
        index_Y_After[4]) );
  ADDHX1 U933 ( .A(n718), .B(\r361/carry[4] ), .CO(\r361/carry[5] ), .S(
        index_X_After[4]) );
  NAND2X1 U934 ( .A(n1092), .B(n1091), .Y(n1095) );
  CLKBUFX3 U935 ( .A(n1112), .Y(n731) );
  AO22XL U936 ( .A0(n1136), .A1(n709), .B0(cdata_rd[19]), .B1(n710), .Y(n377)
         );
  NAND2X1 U937 ( .A(n877), .B(n876), .Y(n383) );
  AOI2BB2X1 U938 ( .B0(N1094), .B1(n727), .A0N(n1033), .A1N(n875), .Y(n876) );
  AOI2BB2X1 U939 ( .B0(N733), .B1(n726), .A0N(n720), .A1N(n874), .Y(n877) );
  AOI2BB2X1 U940 ( .B0(N1104), .B1(n727), .A0N(n722), .A1N(n1017), .Y(n1018)
         );
  AOI2BB2X1 U941 ( .B0(N1103), .B1(n728), .A0N(n722), .A1N(n1020), .Y(n1021)
         );
  NAND2X1 U942 ( .A(n897), .B(n896), .Y(n388) );
  AOI2BB2X1 U943 ( .B0(N1089), .B1(n727), .A0N(n722), .A1N(n895), .Y(n896) );
  AOI2BB2X1 U944 ( .B0(N728), .B1(n726), .A0N(n720), .A1N(n894), .Y(n897) );
  NAND2X1 U945 ( .A(n893), .B(n892), .Y(n387) );
  AOI2BB2X1 U946 ( .B0(N1090), .B1(n727), .A0N(n722), .A1N(n891), .Y(n892) );
  AOI2BB2X1 U947 ( .B0(N729), .B1(n726), .A0N(n720), .A1N(n890), .Y(n893) );
  AOI2BB2X1 U948 ( .B0(N1100), .B1(n727), .A0N(n723), .A1N(n1032), .Y(n1034)
         );
  NAND2X1 U949 ( .A(n873), .B(n872), .Y(n382) );
  AOI2BB2X1 U950 ( .B0(N1095), .B1(n727), .A0N(n723), .A1N(n871), .Y(n872) );
  NAND2X1 U951 ( .A(n885), .B(n884), .Y(n385) );
  AOI2BB2X1 U952 ( .B0(N1092), .B1(n727), .A0N(n722), .A1N(n883), .Y(n884) );
  AOI2BB2X1 U953 ( .B0(N731), .B1(n726), .A0N(n720), .A1N(n882), .Y(n885) );
  NAND2X1 U954 ( .A(n1026), .B(n1025), .Y(n374) );
  AOI2BB2X1 U955 ( .B0(N1102), .B1(n728), .A0N(n722), .A1N(n1024), .Y(n1025)
         );
  NAND2X1 U956 ( .A(n1030), .B(n1029), .Y(n375) );
  AOI2BB2X1 U957 ( .B0(N1101), .B1(n727), .A0N(n722), .A1N(n1028), .Y(n1029)
         );
  NAND2X1 U958 ( .A(n889), .B(n888), .Y(n386) );
  AOI2BB2X1 U959 ( .B0(N1091), .B1(n727), .A0N(n723), .A1N(n887), .Y(n888) );
  AOI2BB2X1 U960 ( .B0(N730), .B1(n726), .A0N(n720), .A1N(n886), .Y(n889) );
  NAND2X1 U961 ( .A(n1005), .B(n1004), .Y(n378) );
  AOI2BB2X1 U962 ( .B0(N1099), .B1(n727), .A0N(n722), .A1N(n1003), .Y(n1004)
         );
  NAND2X1 U963 ( .A(n1001), .B(n1000), .Y(n379) );
  AOI2BB2X1 U964 ( .B0(N1098), .B1(n728), .A0N(n722), .A1N(n999), .Y(n1000) );
  NAND2X1 U965 ( .A(n865), .B(n864), .Y(n380) );
  AOI2BB2X1 U966 ( .B0(N1097), .B1(n727), .A0N(n722), .A1N(n863), .Y(n864) );
  NAND2X1 U967 ( .A(n869), .B(n868), .Y(n381) );
  AOI2BB2X1 U968 ( .B0(N1096), .B1(n727), .A0N(n723), .A1N(n867), .Y(n868) );
  NAND2X1 U969 ( .A(n881), .B(n880), .Y(n384) );
  AOI2BB2X1 U970 ( .B0(N1093), .B1(n727), .A0N(n1033), .A1N(n879), .Y(n880) );
  AOI2BB2X1 U971 ( .B0(N732), .B1(n726), .A0N(n720), .A1N(n878), .Y(n881) );
  NAND2X1 U972 ( .A(convTemp[43]), .B(n1037), .Y(n1038) );
  CLKINVX1 U973 ( .A(n708), .Y(n1108) );
  NAND3BX1 U974 ( .AN(n1051), .B(n262), .C(n696), .Y(n449) );
  NAND2XL U975 ( .A(n1160), .B(n264), .Y(n262) );
  NAND3BX1 U976 ( .AN(counterRead[2]), .B(n1006), .C(n101), .Y(n809) );
  NAND3BX1 U977 ( .AN(n767), .B(n766), .C(n765), .Y(next_State[0]) );
  CLKMX2X2 U978 ( .A(n770), .B(n758), .S0(n682), .Y(n767) );
  AND3X2 U979 ( .A(n1110), .B(n769), .C(n695), .Y(n765) );
  OAI221XL U980 ( .A0(n40), .A1(n1071), .B0(n40), .B1(n1070), .C0(n1069), .Y(
        n424) );
  OA22X1 U981 ( .A0(n708), .A1(n610), .B0(n43), .B1(n1111), .Y(n1069) );
  NAND4X1 U982 ( .A(n269), .B(n1054), .C(n1053), .D(n1052), .Y(n451) );
  NAND2XL U983 ( .A(n1158), .B(n264), .Y(n269) );
  OAI221XL U984 ( .A0(n1111), .A1(n39), .B0(n1109), .B1(n38), .C0(n198), .Y(
        n414) );
  AOI2BB1X1 U985 ( .A0N(n708), .A1N(n642), .B0(n795), .Y(n198) );
  NAND3X1 U986 ( .A(n265), .B(n698), .C(n1107), .Y(n450) );
  CLKINVX1 U987 ( .A(n1051), .Y(n1107) );
  NAND2XL U988 ( .A(n1159), .B(n264), .Y(n265) );
  NAND2X1 U989 ( .A(n937), .B(n936), .Y(n398) );
  AOI2BB2X1 U990 ( .B0(N1079), .B1(n728), .A0N(n722), .A1N(n935), .Y(n936) );
  AOI2BB2X1 U991 ( .B0(N718), .B1(n725), .A0N(n721), .A1N(n934), .Y(n937) );
  NAND2X1 U992 ( .A(n941), .B(n940), .Y(n399) );
  AOI2BB2X1 U993 ( .B0(N1078), .B1(n728), .A0N(n723), .A1N(n939), .Y(n940) );
  AOI2BB2X1 U994 ( .B0(N717), .B1(n725), .A0N(n721), .A1N(n938), .Y(n941) );
  NAND2X1 U995 ( .A(n933), .B(n932), .Y(n397) );
  AOI2BB2X1 U996 ( .B0(N1080), .B1(n728), .A0N(n722), .A1N(n931), .Y(n932) );
  AOI2BB2X1 U997 ( .B0(N719), .B1(n725), .A0N(n721), .A1N(n930), .Y(n933) );
  NAND2X1 U998 ( .A(n913), .B(n912), .Y(n392) );
  AOI2BB2X1 U999 ( .B0(N1085), .B1(n728), .A0N(n723), .A1N(n911), .Y(n912) );
  NAND2X1 U1000 ( .A(n917), .B(n916), .Y(n393) );
  AOI2BB2X1 U1001 ( .B0(N1084), .B1(n728), .A0N(n723), .A1N(n915), .Y(n916) );
  AOI2BB2X1 U1002 ( .B0(N723), .B1(n726), .A0N(n721), .A1N(n914), .Y(n917) );
  NAND2X1 U1003 ( .A(n921), .B(n920), .Y(n394) );
  AOI2BB2X1 U1004 ( .B0(N1083), .B1(n728), .A0N(n723), .A1N(n919), .Y(n920) );
  AOI2BB2X1 U1005 ( .B0(N722), .B1(n726), .A0N(n721), .A1N(n918), .Y(n921) );
  NAND2X1 U1006 ( .A(n909), .B(n908), .Y(n391) );
  AOI2BB2X1 U1007 ( .B0(N1086), .B1(n727), .A0N(n723), .A1N(n907), .Y(n908) );
  NAND2X1 U1008 ( .A(n929), .B(n928), .Y(n396) );
  AOI2BB2X1 U1009 ( .B0(N1081), .B1(n728), .A0N(n1033), .A1N(n927), .Y(n928)
         );
  AOI2BB2X1 U1010 ( .B0(N720), .B1(n725), .A0N(n721), .A1N(n926), .Y(n929) );
  NAND2X1 U1011 ( .A(n901), .B(n900), .Y(n389) );
  AOI2BB2X1 U1012 ( .B0(N1088), .B1(n727), .A0N(n1033), .A1N(n899), .Y(n900)
         );
  NAND2X1 U1013 ( .A(n905), .B(n904), .Y(n390) );
  AOI2BB2X1 U1014 ( .B0(N1087), .B1(n727), .A0N(n1033), .A1N(n903), .Y(n904)
         );
  NAND2X1 U1015 ( .A(n925), .B(n924), .Y(n395) );
  AOI2BB2X1 U1016 ( .B0(N1082), .B1(n728), .A0N(n722), .A1N(n923), .Y(n924) );
  AOI2BB2X1 U1017 ( .B0(N721), .B1(n726), .A0N(n721), .A1N(n922), .Y(n925) );
  NAND2X1 U1018 ( .A(n206), .B(n207), .Y(n420) );
  AOI222XL U1019 ( .A0(n713), .A1(n793), .B0(n142), .B1(N314), .C0(n792), .C1(
        n714), .Y(n207) );
  OA22X1 U1020 ( .A0(n708), .A1(n632), .B0(n791), .B1(n1071), .Y(n206) );
  CLKINVX1 U1021 ( .A(n714), .Y(n791) );
  OAI221XL U1022 ( .A0(n1110), .A1(n38), .B0(n1109), .B1(n37), .C0(n201), .Y(
        n415) );
  OA22X1 U1023 ( .A0(n708), .A1(n620), .B0(n38), .B1(n1071), .Y(n201) );
  OAI221XL U1024 ( .A0(n1110), .A1(n37), .B0(n1109), .B1(n36), .C0(n202), .Y(
        n416) );
  OA22X1 U1025 ( .A0(n708), .A1(n618), .B0(n37), .B1(n1071), .Y(n202) );
  OAI221XL U1026 ( .A0(n1110), .A1(n36), .B0(n1109), .B1(n35), .C0(n203), .Y(
        n417) );
  OA22X1 U1027 ( .A0(n708), .A1(n616), .B0(n794), .B1(n1071), .Y(n203) );
  CLKINVX1 U1028 ( .A(n717), .Y(n794) );
  OAI221XL U1029 ( .A0(n1110), .A1(n35), .B0(n1109), .B1(n28), .C0(n204), .Y(
        n418) );
  OA22X1 U1030 ( .A0(n708), .A1(n614), .B0(n35), .B1(n1071), .Y(n204) );
  OAI221XL U1031 ( .A0(n1110), .A1(n28), .B0(n1109), .B1(n46), .C0(n205), .Y(
        n419) );
  OA22X1 U1032 ( .A0(n708), .A1(n612), .B0(n28), .B1(n1071), .Y(n205) );
  NAND2X1 U1033 ( .A(n945), .B(n944), .Y(n400) );
  AOI2BB2X1 U1034 ( .B0(N1077), .B1(n728), .A0N(n723), .A1N(n943), .Y(n944) );
  AOI2BB2X1 U1035 ( .B0(N716), .B1(n725), .A0N(n721), .A1N(n942), .Y(n945) );
  NAND2X1 U1036 ( .A(n949), .B(n948), .Y(n401) );
  AOI2BB2X1 U1037 ( .B0(N1076), .B1(n728), .A0N(n723), .A1N(n947), .Y(n948) );
  AOI2BB2X1 U1038 ( .B0(N715), .B1(n725), .A0N(n721), .A1N(n946), .Y(n949) );
  NAND2X1 U1039 ( .A(n961), .B(n960), .Y(n404) );
  AOI2BB2X1 U1040 ( .B0(N1073), .B1(n686), .A0N(n723), .A1N(n959), .Y(n960) );
  AOI2BB2X1 U1041 ( .B0(N712), .B1(n725), .A0N(n1031), .A1N(n958), .Y(n961) );
  CLKINVX1 U1042 ( .A(reset), .Y(n1112) );
  NAND2X1 U1043 ( .A(n953), .B(n952), .Y(n402) );
  AOI2BB2X1 U1044 ( .B0(N1075), .B1(n728), .A0N(n723), .A1N(n951), .Y(n952) );
  AOI2BB2X1 U1045 ( .B0(N714), .B1(n725), .A0N(n721), .A1N(n950), .Y(n953) );
  NAND2X1 U1046 ( .A(n957), .B(n956), .Y(n403) );
  AOI2BB2X1 U1047 ( .B0(N1074), .B1(n728), .A0N(n723), .A1N(n955), .Y(n956) );
  AOI2BB2X1 U1048 ( .B0(N713), .B1(n725), .A0N(n721), .A1N(n954), .Y(n957) );
  NAND3BX1 U1049 ( .AN(current_State[1]), .B(n81), .C(n693), .Y(n787) );
  NAND2X1 U1050 ( .A(n965), .B(n964), .Y(n405) );
  AOI2BB2X1 U1051 ( .B0(N1072), .B1(n686), .A0N(n723), .A1N(n963), .Y(n964) );
  AOI2BB2X1 U1052 ( .B0(N711), .B1(n725), .A0N(n1031), .A1N(n962), .Y(n965) );
  NAND2X1 U1053 ( .A(n973), .B(n972), .Y(n407) );
  AOI2BB2X1 U1054 ( .B0(N1070), .B1(n686), .A0N(n723), .A1N(n971), .Y(n972) );
  AOI2BB2X1 U1055 ( .B0(N709), .B1(n724), .A0N(n1031), .A1N(n970), .Y(n973) );
  AO21XL U1056 ( .A0(n1132), .A1(n1105), .B0(ready), .Y(n452) );
  NAND2X1 U1057 ( .A(n969), .B(n968), .Y(n406) );
  AOI2BB2X1 U1058 ( .B0(N1071), .B1(n686), .A0N(n723), .A1N(n967), .Y(n968) );
  AOI2BB2X1 U1059 ( .B0(N710), .B1(n725), .A0N(n720), .A1N(n966), .Y(n969) );
  NAND2X1 U1060 ( .A(n977), .B(n976), .Y(n408) );
  AOI2BB2X1 U1061 ( .B0(N1069), .B1(n686), .A0N(n723), .A1N(n975), .Y(n976) );
  AOI2BB2X1 U1062 ( .B0(N708), .B1(n724), .A0N(n721), .A1N(n974), .Y(n977) );
  NAND2X1 U1063 ( .A(n981), .B(n980), .Y(n409) );
  AOI2BB2X1 U1064 ( .B0(N1068), .B1(n686), .A0N(n723), .A1N(n979), .Y(n980) );
  AOI2BB2X1 U1065 ( .B0(N707), .B1(n724), .A0N(n721), .A1N(n978), .Y(n981) );
  BUFX4 U1066 ( .A(n120), .Y(n711) );
  NOR2X1 U1067 ( .A(roundTemp[20]), .B(n1111), .Y(n120) );
  NAND2X1 U1068 ( .A(n80), .B(n1009), .Y(n1070) );
  NAND4X1 U1069 ( .A(n775), .B(n774), .C(n773), .D(n772), .Y(next_State[1]) );
  OA22X1 U1070 ( .A0(n351), .A1(n788), .B0(n1124), .B1(n787), .Y(n772) );
  NAND3BX1 U1071 ( .AN(N314), .B(n359), .C(n783), .Y(n763) );
  NAND4X1 U1072 ( .A(n718), .B(n717), .C(N559), .D(n367), .Y(n294) );
  NOR3X1 U1073 ( .A(n37), .B(N279), .C(n38), .Y(n367) );
  NAND2X1 U1074 ( .A(n985), .B(n984), .Y(n410) );
  AOI2BB2X1 U1075 ( .B0(N1067), .B1(n686), .A0N(n723), .A1N(n983), .Y(n984) );
  AOI2BB2X1 U1076 ( .B0(N706), .B1(n724), .A0N(n720), .A1N(n982), .Y(n985) );
  NAND2X1 U1077 ( .A(n989), .B(n988), .Y(n411) );
  AOI2BB2X1 U1078 ( .B0(N1066), .B1(n686), .A0N(n723), .A1N(n987), .Y(n988) );
  AOI2BB2X1 U1079 ( .B0(N705), .B1(n724), .A0N(n721), .A1N(n986), .Y(n989) );
  NAND2X1 U1080 ( .A(n993), .B(n992), .Y(n412) );
  AOI2BB2X1 U1081 ( .B0(N1065), .B1(n686), .A0N(n723), .A1N(n991), .Y(n992) );
  AOI2BB2X1 U1082 ( .B0(N704), .B1(n724), .A0N(n1031), .A1N(n990), .Y(n993) );
  NAND2X1 U1083 ( .A(n997), .B(n996), .Y(n413) );
  AOI2BB2X1 U1084 ( .B0(N1064), .B1(n686), .A0N(n722), .A1N(n995), .Y(n996) );
  AOI2BB2X1 U1085 ( .B0(N703), .B1(n724), .A0N(n720), .A1N(n994), .Y(n997) );
  NAND3BX1 U1086 ( .AN(n78), .B(n81), .C(n704), .Y(n1065) );
  MXI2X1 U1087 ( .A(n634), .B(n1104), .S0(n706), .Y(n448) );
  AOI222XL U1088 ( .A0(index_Y_Before[5]), .A1(n1102), .B0(n716), .B1(n1101), 
        .C0(index_Y_After[5]), .C1(n561), .Y(n1104) );
  MXI2X1 U1089 ( .A(n584), .B(n1096), .S0(n706), .Y(n444) );
  AOI222XL U1090 ( .A0(index_Y_Before[1]), .A1(n1102), .B0(n714), .B1(n1101), 
        .C0(index_Y_After[1]), .C1(n561), .Y(n1096) );
  MXI2X1 U1091 ( .A(n582), .B(n1097), .S0(n706), .Y(n445) );
  AOI222XL U1092 ( .A0(index_Y_Before[2]), .A1(n1102), .B0(n713), .B1(n1101), 
        .C0(index_Y_After[2]), .C1(n561), .Y(n1097) );
  MXI2X1 U1093 ( .A(n636), .B(n1099), .S0(n706), .Y(n447) );
  AOI222XL U1094 ( .A0(index_Y_Before[4]), .A1(n1102), .B0(n715), .B1(n1101), 
        .C0(index_Y_After[4]), .C1(n561), .Y(n1099) );
  NAND3BX1 U1095 ( .AN(n78), .B(n79), .C(n701), .Y(n1066) );
  CLKINVX1 U1096 ( .A(n755), .Y(n756) );
  OAI21XL U1097 ( .A0(n28), .A1(n277), .B0(n293), .Y(n463) );
  AOI22X1 U1098 ( .A0(n279), .A1(index_X_After[5]), .B0(N284), .B1(n697), .Y(
        n293) );
  OAI21XL U1099 ( .A0(n40), .A1(n285), .B0(n296), .Y(n464) );
  AOI22X1 U1100 ( .A0(n287), .A1(index_Y_After[5]), .B0(N319), .B1(n473), .Y(
        n296) );
  NAND3X1 U1101 ( .A(n46), .B(n45), .C(n47), .Y(n192) );
  NOR2BX1 U1102 ( .AN(n359), .B(n47), .Y(n185) );
  NAND4X1 U1103 ( .A(N556), .B(N555), .C(n717), .D(n360), .Y(n191) );
  NOR3X1 U1104 ( .A(n39), .B(n35), .C(n28), .Y(n360) );
  NAND4X1 U1105 ( .A(n38), .B(n37), .C(n39), .D(n194), .Y(n184) );
  NOR3X1 U1106 ( .A(n717), .B(N559), .C(n718), .Y(n194) );
  MXI2X1 U1107 ( .A(n638), .B(n1090), .S0(n706), .Y(n442) );
  AOI222XL U1108 ( .A0(index_X_Before[5]), .A1(n1089), .B0(N559), .B1(n1088), 
        .C0(index_X_After[5]), .C1(n1087), .Y(n1090) );
  OAI21XL U1109 ( .A0(n36), .A1(n277), .B0(n281), .Y(n454) );
  AOI22X1 U1110 ( .A0(n279), .A1(index_X_After[3]), .B0(N282), .B1(n697), .Y(
        n281) );
  OAI21XL U1111 ( .A0(n35), .A1(n277), .B0(n278), .Y(n453) );
  AOI22X1 U1112 ( .A0(n279), .A1(index_X_After[4]), .B0(N283), .B1(n697), .Y(
        n278) );
  MXI2X1 U1113 ( .A(n588), .B(n1083), .S0(n706), .Y(n438) );
  AOI222XL U1114 ( .A0(index_X_Before[1]), .A1(n1089), .B0(N555), .B1(n1088), 
        .C0(index_X_After[1]), .C1(n1087), .Y(n1083) );
  MXI2X1 U1115 ( .A(n586), .B(n1084), .S0(n706), .Y(n439) );
  AOI222XL U1116 ( .A0(index_X_Before[2]), .A1(n1089), .B0(N556), .B1(n1088), 
        .C0(index_X_After[2]), .C1(n1087), .Y(n1084) );
  MXI2X1 U1117 ( .A(n624), .B(n1085), .S0(n706), .Y(n440) );
  AOI222XL U1118 ( .A0(index_X_Before[3]), .A1(n1089), .B0(n717), .B1(n1088), 
        .C0(index_X_After[3]), .C1(n1087), .Y(n1085) );
  MXI2X1 U1119 ( .A(n640), .B(n1086), .S0(n706), .Y(n441) );
  AOI222XL U1120 ( .A0(index_X_Before[4]), .A1(n1089), .B0(n718), .B1(n1088), 
        .C0(index_X_After[4]), .C1(n1087), .Y(n1086) );
  MXI2X1 U1121 ( .A(n622), .B(n1098), .S0(n706), .Y(n446) );
  AOI222XL U1122 ( .A0(index_Y_Before[3]), .A1(n1102), .B0(n712), .B1(n1101), 
        .C0(index_Y_After[3]), .C1(n561), .Y(n1098) );
  OAI21XL U1123 ( .A0(n37), .A1(n277), .B0(n282), .Y(n455) );
  AOI22X1 U1124 ( .A0(n279), .A1(index_X_After[2]), .B0(N281), .B1(n697), .Y(
        n282) );
  OAI21XL U1125 ( .A0(n38), .A1(n277), .B0(n283), .Y(n456) );
  AOI22X1 U1126 ( .A0(n279), .A1(index_X_After[1]), .B0(n38), .B1(n697), .Y(
        n283) );
  OAI21XL U1127 ( .A0(n39), .A1(n277), .B0(n284), .Y(n457) );
  AOI22X1 U1128 ( .A0(n279), .A1(n39), .B0(N279), .B1(n697), .Y(n284) );
  OAI21XL U1129 ( .A0(n44), .A1(n285), .B0(n289), .Y(n459) );
  AOI22X1 U1130 ( .A0(n287), .A1(index_Y_After[3]), .B0(N317), .B1(n473), .Y(
        n289) );
  OAI21XL U1131 ( .A0(n45), .A1(n285), .B0(n290), .Y(n460) );
  AOI22X1 U1132 ( .A0(n287), .A1(index_Y_After[2]), .B0(N316), .B1(n473), .Y(
        n290) );
  OAI21XL U1133 ( .A0(n46), .A1(n285), .B0(n291), .Y(n461) );
  AOI22X1 U1134 ( .A0(n287), .A1(index_Y_After[1]), .B0(n791), .B1(n473), .Y(
        n291) );
  OAI21XL U1135 ( .A0(n47), .A1(n285), .B0(n292), .Y(n462) );
  AOI22X1 U1136 ( .A0(n287), .A1(n47), .B0(N314), .B1(n473), .Y(n292) );
  OAI21XL U1137 ( .A0(n43), .A1(n285), .B0(n286), .Y(n458) );
  AOI22X1 U1138 ( .A0(n287), .A1(index_Y_After[4]), .B0(N318), .B1(n473), .Y(
        n286) );
  MX2XL U1139 ( .A(n1134), .B(n1082), .S0(n706), .Y(n437) );
  CLKMX2X2 U1140 ( .A(n1081), .B(n1088), .S0(N279), .Y(n1082) );
  NAND2X1 U1141 ( .A(n1078), .B(n1077), .Y(n1081) );
  CLKINVX1 U1142 ( .A(n1089), .Y(n1077) );
  AND4X1 U1143 ( .A(n716), .B(n715), .C(n368), .D(n712), .Y(n359) );
  NOR2X1 U1144 ( .A(n46), .B(n45), .Y(n368) );
  MXI2X1 U1145 ( .A(n702), .B(n703), .S0(n706), .Y(n443) );
  CLKBUFX3 U1146 ( .A(N562), .Y(n712) );
  CLKBUFX3 U1147 ( .A(N563), .Y(n715) );
  CLKBUFX3 U1148 ( .A(N557), .Y(n717) );
  CLKBUFX3 U1149 ( .A(N558), .Y(n718) );
  CLKBUFX3 U1150 ( .A(N560), .Y(n714) );
  CLKBUFX3 U1151 ( .A(N564), .Y(n716) );
  NAND2X1 U1152 ( .A(n689), .B(n101), .Y(n1047) );
  NAND2X1 U1153 ( .A(n689), .B(n99), .Y(n1062) );
  OAI221XL U1154 ( .A0(N279), .A1(n1048), .B0(n39), .B1(n1047), .C0(n1041), 
        .Y(n425) );
  OA22X1 U1155 ( .A0(n38), .A1(n472), .B0(n1060), .B1(n608), .Y(n1041) );
  OAI221XL U1156 ( .A0(n1129), .A1(n1048), .B0(n38), .B1(n1047), .C0(n1042), 
        .Y(n426) );
  CLKINVX1 U1157 ( .A(index_X_After[1]), .Y(n1129) );
  OA22X1 U1158 ( .A0(n37), .A1(n472), .B0(n1060), .B1(n606), .Y(n1042) );
  OAI221XL U1159 ( .A0(n1128), .A1(n1048), .B0(n37), .B1(n1047), .C0(n1043), 
        .Y(n427) );
  CLKINVX1 U1160 ( .A(index_X_After[2]), .Y(n1128) );
  OA22X1 U1161 ( .A0(n36), .A1(n472), .B0(n1060), .B1(n604), .Y(n1043) );
  OAI221XL U1162 ( .A0(n1127), .A1(n1048), .B0(n36), .B1(n1047), .C0(n1044), 
        .Y(n428) );
  CLKINVX1 U1163 ( .A(index_X_After[3]), .Y(n1127) );
  OA22X1 U1164 ( .A0(n35), .A1(n472), .B0(n1060), .B1(n602), .Y(n1044) );
  OAI221XL U1165 ( .A0(n1126), .A1(n1048), .B0(n35), .B1(n1047), .C0(n1045), 
        .Y(n429) );
  CLKINVX1 U1166 ( .A(index_X_After[4]), .Y(n1126) );
  OA22X1 U1167 ( .A0(n28), .A1(n472), .B0(n1060), .B1(n600), .Y(n1045) );
  OAI221XL U1168 ( .A0(n1125), .A1(n1048), .B0(n28), .B1(n1047), .C0(n1046), 
        .Y(n430) );
  CLKINVX1 U1169 ( .A(index_X_After[5]), .Y(n1125) );
  OA22X1 U1170 ( .A0(n46), .A1(n472), .B0(n1060), .B1(n598), .Y(n1046) );
  OAI221XL U1171 ( .A0(N314), .A1(n1063), .B0(n47), .B1(n1062), .C0(n1055), 
        .Y(n431) );
  OA22X1 U1172 ( .A0(n45), .A1(n472), .B0(n1060), .B1(n596), .Y(n1055) );
  OAI221XL U1173 ( .A0(n1057), .A1(n1063), .B0(n46), .B1(n1062), .C0(n1056), 
        .Y(n432) );
  CLKINVX1 U1174 ( .A(index_Y_After[1]), .Y(n1057) );
  OA22X1 U1175 ( .A0(n44), .A1(n472), .B0(n1060), .B1(n594), .Y(n1056) );
  OAI221XL U1176 ( .A0(n1059), .A1(n1063), .B0(n45), .B1(n1062), .C0(n1058), 
        .Y(n433) );
  CLKINVX1 U1177 ( .A(index_Y_After[2]), .Y(n1059) );
  OA22X1 U1178 ( .A0(n43), .A1(n472), .B0(n1060), .B1(n592), .Y(n1058) );
  OAI221XL U1179 ( .A0(n1064), .A1(n1063), .B0(n44), .B1(n1062), .C0(n1061), 
        .Y(n434) );
  CLKINVX1 U1180 ( .A(index_Y_After[3]), .Y(n1064) );
  OA22X1 U1181 ( .A0(n40), .A1(n472), .B0(n1060), .B1(n590), .Y(n1061) );
  OAI221XL U1182 ( .A0(n1131), .A1(n1063), .B0(n43), .B1(n1062), .C0(n235), 
        .Y(n435) );
  CLKINVX1 U1183 ( .A(index_Y_After[4]), .Y(n1131) );
  NAND2XL U1184 ( .A(n1157), .B(n1106), .Y(n235) );
  OAI221XL U1185 ( .A0(n1130), .A1(n1063), .B0(n40), .B1(n1062), .C0(n236), 
        .Y(n436) );
  CLKINVX1 U1186 ( .A(index_Y_After[5]), .Y(n1130) );
  NAND2XL U1187 ( .A(n1156), .B(n1106), .Y(n236) );
  ADDHX1 U1188 ( .A(n714), .B(N314), .CO(\r363/carry[2] ), .S(index_Y_After[1]) );
  ADDHX1 U1189 ( .A(N555), .B(N279), .CO(\r361/carry[2] ), .S(index_X_After[1]) );
  ADDHX1 U1190 ( .A(N556), .B(\r361/carry[2] ), .CO(\r361/carry[3] ), .S(
        index_X_After[2]) );
  CLKBUFX3 U1191 ( .A(N561), .Y(n713) );
  NAND2X2 U1192 ( .A(n787), .B(n788), .Y(n142) );
  NAND2X2 U1193 ( .A(n1076), .B(n559), .Y(n1101) );
  XOR2X1 U1194 ( .A(n716), .B(\add_153_S2/carry[5] ), .Y(N319) );
  AND2X1 U1195 ( .A(\add_153_S2/carry[4] ), .B(n715), .Y(\add_153_S2/carry[5] ) );
  XOR2X1 U1196 ( .A(n715), .B(\add_153_S2/carry[4] ), .Y(N318) );
  AND2X1 U1197 ( .A(\add_153_S2/carry[3] ), .B(n712), .Y(\add_153_S2/carry[4] ) );
  XOR2X1 U1198 ( .A(n712), .B(\add_153_S2/carry[3] ), .Y(N317) );
  AND2X1 U1199 ( .A(n714), .B(n713), .Y(\add_153_S2/carry[3] ) );
  XOR2X1 U1200 ( .A(n713), .B(n714), .Y(N316) );
  XOR2X1 U1201 ( .A(N559), .B(\add_140/carry[5] ), .Y(N284) );
  AND2X1 U1202 ( .A(\add_140/carry[4] ), .B(n718), .Y(\add_140/carry[5] ) );
  XOR2X1 U1203 ( .A(n718), .B(\add_140/carry[4] ), .Y(N283) );
  AND2X1 U1204 ( .A(\add_140/carry[3] ), .B(n717), .Y(\add_140/carry[4] ) );
  XOR2X1 U1205 ( .A(n717), .B(\add_140/carry[3] ), .Y(N282) );
  AND2X1 U1206 ( .A(N555), .B(N556), .Y(\add_140/carry[3] ) );
  XOR2X1 U1207 ( .A(N556), .B(N555), .Y(N281) );
  XOR2X1 U1208 ( .A(\r361/carry[5] ), .B(N559), .Y(index_X_After[5]) );
  XOR2X1 U1209 ( .A(\r363/carry[5] ), .B(n716), .Y(index_Y_After[5]) );
  NAND2BX1 U1210 ( .AN(N555), .B(n39), .Y(n1114) );
  OAI2BB1X1 U1211 ( .A0N(N279), .A1N(N555), .B0(n1114), .Y(index_X_Before[1])
         );
  NOR2X1 U1212 ( .A(n1114), .B(N556), .Y(n1115) );
  AO21X1 U1213 ( .A0(n1114), .A1(N556), .B0(n1115), .Y(index_X_Before[2]) );
  NAND2X1 U1214 ( .A(n1115), .B(n36), .Y(n1116) );
  OAI21XL U1215 ( .A0(n1115), .A1(n794), .B0(n1116), .Y(index_X_Before[3]) );
  XNOR2X1 U1216 ( .A(n718), .B(n1116), .Y(index_X_Before[4]) );
  NOR2X1 U1217 ( .A(n718), .B(n1116), .Y(n1117) );
  XOR2X1 U1218 ( .A(N559), .B(n1117), .Y(index_X_Before[5]) );
  NAND2BX1 U1219 ( .AN(n714), .B(n47), .Y(n1118) );
  OAI2BB1X1 U1220 ( .A0N(N314), .A1N(n714), .B0(n1118), .Y(index_Y_Before[1])
         );
  NOR2X1 U1221 ( .A(n1118), .B(n713), .Y(n1119) );
  AO21X1 U1222 ( .A0(n1118), .A1(n713), .B0(n1119), .Y(index_Y_Before[2]) );
  NAND2X1 U1223 ( .A(n1119), .B(n44), .Y(n1120) );
  OAI21XL U1224 ( .A0(n1119), .A1(n44), .B0(n1120), .Y(index_Y_Before[3]) );
  XNOR2X1 U1225 ( .A(n715), .B(n1120), .Y(index_Y_Before[4]) );
  NOR2X1 U1226 ( .A(n715), .B(n1120), .Y(n1121) );
  XOR2X1 U1227 ( .A(n716), .B(n1121), .Y(index_Y_Before[5]) );
  CONV_DW01_add_0 add_395 ( .A(convTemp), .B({1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, n707, n707, n707, n707, 1'b0, n707, n707, 1'b1, 1'b0, 
        1'b0, 1'b1, n1123, n707, 1'b0, 1'b0, 1'b1, 1'b0, n707, 1'b0, n707, 
        1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 1'b0, 
        1'b0, 1'b0, 1'b0, 1'b0}), .CI(1'b0), .SUM({N1107, N1106, N1105, N1104, 
        N1103, N1102, N1101, N1100, N1099, N1098, N1097, N1096, N1095, N1094, 
        N1093, N1092, N1091, N1090, N1089, N1088, N1087, N1086, N1085, N1084, 
        N1083, N1082, N1081, N1080, N1079, N1078, N1077, N1076, N1075, N1074, 
        N1073, N1072, N1071, N1070, N1069, N1068, N1067, N1066, N1065, N1064})
         );
  CONV_DW_cmp_0 gt_363 ( .A(cdata_rd), .B({n1136, n1137, n1138, n1139, n1140, 
        n1141, n1142, n1143, n1144, n1145, n1146, n1147, n1148, n1149, n1150, 
        n1151, n1152, n1153, n1154, n1155}), .TC(1'b0), .GE_LT(1'b0), 
        .GE_GT_EQ(1'b1), .GE_LT_GT_LE(N610) );
  CONV_DW01_inc_1 add_38 ( .A(convTemp[35:15]), .SUM({roundTemp, 
        SYNOPSYS_UNCONNECTED__0}) );
  CONV_DW_mult_tc_2 mult_375 ( .a({kernelTemp[19], kernelTemp[19], 
        kernelTemp[19], kernelTemp[19], kernelTemp[15:0]}), .b(idataTemp), 
        .product({mulTemp_43, mulTemp}) );
  CONV_DW01_add_5 r370 ( .A(convTemp), .B({mulTemp_43, mulTemp_43, mulTemp_43, 
        mulTemp_43, mulTemp_43, mulTemp[38:29], n560, mulTemp[27:16], n558, 
        mulTemp[14:7], n557, mulTemp[5:0]}), .CI(1'b0), .SUM({N746, N745, N744, 
        N743, N742, N741, N740, N739, N738, N737, N736, N735, N734, N733, N732, 
        N731, N730, N729, N728, N727, N726, N725, N724, N723, N722, N721, N720, 
        N719, N718, N717, N716, N715, N714, N713, N712, N711, N710, N709, N708, 
        N707, N706, N705, N704, N703}) );
  DFFRX1 crd_reg ( .D(N430), .CK(clk), .RN(n1112), .QN(n500) );
  DFFRX1 \iaddr_reg[7]  ( .D(n444), .CK(clk), .RN(n1112), .Q(n1163), .QN(n584)
         );
  INVXL U545 ( .A(n1163), .Y(n1161) );
  INVX12 U638 ( .A(n1161), .Y(iaddr[7]) );
endmodule

